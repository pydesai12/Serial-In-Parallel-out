
module serial_DW01_inc_3 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  CHA1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CHA1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CHA1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CHA1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CHA1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CEOX1 U1 ( .A(carry[6]), .B(A[6]), .Z(SUM[6]) );
  CIVX1 U2 ( .A(A[0]), .Z(SUM[0]) );
endmodule


module serial ( clk, rst, pushin, lastin, datain, pullout, stopout, dataout, 
        lenout );
  output [63:0] dataout;
  output [6:0] lenout;
  input clk, rst, pushin, lastin, datain, pullout;
  output stopout;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N38, N39, N40, N41, N42, \memory[31][70] , \memory[31][69] ,
         \memory[31][68] , \memory[31][67] , \memory[31][66] ,
         \memory[31][65] , \memory[31][64] , \memory[31][63] ,
         \memory[31][62] , \memory[31][61] , \memory[31][60] ,
         \memory[31][59] , \memory[31][58] , \memory[31][57] ,
         \memory[31][56] , \memory[31][55] , \memory[31][54] ,
         \memory[31][53] , \memory[31][52] , \memory[31][51] ,
         \memory[31][50] , \memory[31][49] , \memory[31][48] ,
         \memory[31][47] , \memory[31][46] , \memory[31][45] ,
         \memory[31][44] , \memory[31][43] , \memory[31][42] ,
         \memory[31][41] , \memory[31][40] , \memory[31][39] ,
         \memory[31][38] , \memory[31][37] , \memory[31][36] ,
         \memory[31][35] , \memory[31][34] , \memory[31][33] ,
         \memory[31][32] , \memory[31][31] , \memory[31][30] ,
         \memory[31][29] , \memory[31][28] , \memory[31][27] ,
         \memory[31][26] , \memory[31][25] , \memory[31][24] ,
         \memory[31][23] , \memory[31][22] , \memory[31][21] ,
         \memory[31][20] , \memory[31][19] , \memory[31][18] ,
         \memory[31][17] , \memory[31][16] , \memory[31][15] ,
         \memory[31][14] , \memory[31][13] , \memory[31][12] ,
         \memory[31][11] , \memory[31][10] , \memory[31][9] , \memory[31][8] ,
         \memory[31][7] , \memory[31][6] , \memory[31][5] , \memory[31][4] ,
         \memory[31][3] , \memory[31][2] , \memory[31][1] , \memory[31][0] ,
         \memory[30][70] , \memory[30][69] , \memory[30][68] ,
         \memory[30][67] , \memory[30][66] , \memory[30][65] ,
         \memory[30][64] , \memory[30][63] , \memory[30][62] ,
         \memory[30][61] , \memory[30][60] , \memory[30][59] ,
         \memory[30][58] , \memory[30][57] , \memory[30][56] ,
         \memory[30][55] , \memory[30][54] , \memory[30][53] ,
         \memory[30][52] , \memory[30][51] , \memory[30][50] ,
         \memory[30][49] , \memory[30][48] , \memory[30][47] ,
         \memory[30][46] , \memory[30][45] , \memory[30][44] ,
         \memory[30][43] , \memory[30][42] , \memory[30][41] ,
         \memory[30][40] , \memory[30][39] , \memory[30][38] ,
         \memory[30][37] , \memory[30][36] , \memory[30][35] ,
         \memory[30][34] , \memory[30][33] , \memory[30][32] ,
         \memory[30][31] , \memory[30][30] , \memory[30][29] ,
         \memory[30][28] , \memory[30][27] , \memory[30][26] ,
         \memory[30][25] , \memory[30][24] , \memory[30][23] ,
         \memory[30][22] , \memory[30][21] , \memory[30][20] ,
         \memory[30][19] , \memory[30][18] , \memory[30][17] ,
         \memory[30][16] , \memory[30][15] , \memory[30][14] ,
         \memory[30][13] , \memory[30][12] , \memory[30][11] ,
         \memory[30][10] , \memory[30][9] , \memory[30][8] , \memory[30][7] ,
         \memory[30][6] , \memory[30][5] , \memory[30][4] , \memory[30][3] ,
         \memory[30][2] , \memory[30][1] , \memory[30][0] , \memory[29][70] ,
         \memory[29][69] , \memory[29][68] , \memory[29][67] ,
         \memory[29][66] , \memory[29][65] , \memory[29][64] ,
         \memory[29][63] , \memory[29][62] , \memory[29][61] ,
         \memory[29][60] , \memory[29][59] , \memory[29][58] ,
         \memory[29][57] , \memory[29][56] , \memory[29][55] ,
         \memory[29][54] , \memory[29][53] , \memory[29][52] ,
         \memory[29][51] , \memory[29][50] , \memory[29][49] ,
         \memory[29][48] , \memory[29][47] , \memory[29][46] ,
         \memory[29][45] , \memory[29][44] , \memory[29][43] ,
         \memory[29][42] , \memory[29][41] , \memory[29][40] ,
         \memory[29][39] , \memory[29][38] , \memory[29][37] ,
         \memory[29][36] , \memory[29][35] , \memory[29][34] ,
         \memory[29][33] , \memory[29][32] , \memory[29][31] ,
         \memory[29][30] , \memory[29][29] , \memory[29][28] ,
         \memory[29][27] , \memory[29][26] , \memory[29][25] ,
         \memory[29][24] , \memory[29][23] , \memory[29][22] ,
         \memory[29][21] , \memory[29][20] , \memory[29][19] ,
         \memory[29][18] , \memory[29][17] , \memory[29][16] ,
         \memory[29][15] , \memory[29][14] , \memory[29][13] ,
         \memory[29][12] , \memory[29][11] , \memory[29][10] , \memory[29][9] ,
         \memory[29][8] , \memory[29][7] , \memory[29][6] , \memory[29][5] ,
         \memory[29][4] , \memory[29][3] , \memory[29][2] , \memory[29][1] ,
         \memory[29][0] , \memory[28][70] , \memory[28][69] , \memory[28][68] ,
         \memory[28][67] , \memory[28][66] , \memory[28][65] ,
         \memory[28][64] , \memory[28][63] , \memory[28][62] ,
         \memory[28][61] , \memory[28][60] , \memory[28][59] ,
         \memory[28][58] , \memory[28][57] , \memory[28][56] ,
         \memory[28][55] , \memory[28][54] , \memory[28][53] ,
         \memory[28][52] , \memory[28][51] , \memory[28][50] ,
         \memory[28][49] , \memory[28][48] , \memory[28][47] ,
         \memory[28][46] , \memory[28][45] , \memory[28][44] ,
         \memory[28][43] , \memory[28][42] , \memory[28][41] ,
         \memory[28][40] , \memory[28][39] , \memory[28][38] ,
         \memory[28][37] , \memory[28][36] , \memory[28][35] ,
         \memory[28][34] , \memory[28][33] , \memory[28][32] ,
         \memory[28][31] , \memory[28][30] , \memory[28][29] ,
         \memory[28][28] , \memory[28][27] , \memory[28][26] ,
         \memory[28][25] , \memory[28][24] , \memory[28][23] ,
         \memory[28][22] , \memory[28][21] , \memory[28][20] ,
         \memory[28][19] , \memory[28][18] , \memory[28][17] ,
         \memory[28][16] , \memory[28][15] , \memory[28][14] ,
         \memory[28][13] , \memory[28][12] , \memory[28][11] ,
         \memory[28][10] , \memory[28][9] , \memory[28][8] , \memory[28][7] ,
         \memory[28][6] , \memory[28][5] , \memory[28][4] , \memory[28][3] ,
         \memory[28][2] , \memory[28][1] , \memory[28][0] , \memory[27][70] ,
         \memory[27][69] , \memory[27][68] , \memory[27][67] ,
         \memory[27][66] , \memory[27][65] , \memory[27][64] ,
         \memory[27][63] , \memory[27][62] , \memory[27][61] ,
         \memory[27][60] , \memory[27][59] , \memory[27][58] ,
         \memory[27][57] , \memory[27][56] , \memory[27][55] ,
         \memory[27][54] , \memory[27][53] , \memory[27][52] ,
         \memory[27][51] , \memory[27][50] , \memory[27][49] ,
         \memory[27][48] , \memory[27][47] , \memory[27][46] ,
         \memory[27][45] , \memory[27][44] , \memory[27][43] ,
         \memory[27][42] , \memory[27][41] , \memory[27][40] ,
         \memory[27][39] , \memory[27][38] , \memory[27][37] ,
         \memory[27][36] , \memory[27][35] , \memory[27][34] ,
         \memory[27][33] , \memory[27][32] , \memory[27][31] ,
         \memory[27][30] , \memory[27][29] , \memory[27][28] ,
         \memory[27][27] , \memory[27][26] , \memory[27][25] ,
         \memory[27][24] , \memory[27][23] , \memory[27][22] ,
         \memory[27][21] , \memory[27][20] , \memory[27][19] ,
         \memory[27][18] , \memory[27][17] , \memory[27][16] ,
         \memory[27][15] , \memory[27][14] , \memory[27][13] ,
         \memory[27][12] , \memory[27][11] , \memory[27][10] , \memory[27][9] ,
         \memory[27][8] , \memory[27][7] , \memory[27][6] , \memory[27][5] ,
         \memory[27][4] , \memory[27][3] , \memory[27][2] , \memory[27][1] ,
         \memory[27][0] , \memory[26][70] , \memory[26][69] , \memory[26][68] ,
         \memory[26][67] , \memory[26][66] , \memory[26][65] ,
         \memory[26][64] , \memory[26][63] , \memory[26][62] ,
         \memory[26][61] , \memory[26][60] , \memory[26][59] ,
         \memory[26][58] , \memory[26][57] , \memory[26][56] ,
         \memory[26][55] , \memory[26][54] , \memory[26][53] ,
         \memory[26][52] , \memory[26][51] , \memory[26][50] ,
         \memory[26][49] , \memory[26][48] , \memory[26][47] ,
         \memory[26][46] , \memory[26][45] , \memory[26][44] ,
         \memory[26][43] , \memory[26][42] , \memory[26][41] ,
         \memory[26][40] , \memory[26][39] , \memory[26][38] ,
         \memory[26][37] , \memory[26][36] , \memory[26][35] ,
         \memory[26][34] , \memory[26][33] , \memory[26][32] ,
         \memory[26][31] , \memory[26][30] , \memory[26][29] ,
         \memory[26][28] , \memory[26][27] , \memory[26][26] ,
         \memory[26][25] , \memory[26][24] , \memory[26][23] ,
         \memory[26][22] , \memory[26][21] , \memory[26][20] ,
         \memory[26][19] , \memory[26][18] , \memory[26][17] ,
         \memory[26][16] , \memory[26][15] , \memory[26][14] ,
         \memory[26][13] , \memory[26][12] , \memory[26][11] ,
         \memory[26][10] , \memory[26][9] , \memory[26][8] , \memory[26][7] ,
         \memory[26][6] , \memory[26][5] , \memory[26][4] , \memory[26][3] ,
         \memory[26][2] , \memory[26][1] , \memory[26][0] , \memory[25][70] ,
         \memory[25][69] , \memory[25][68] , \memory[25][67] ,
         \memory[25][66] , \memory[25][65] , \memory[25][64] ,
         \memory[25][63] , \memory[25][62] , \memory[25][61] ,
         \memory[25][60] , \memory[25][59] , \memory[25][58] ,
         \memory[25][57] , \memory[25][56] , \memory[25][55] ,
         \memory[25][54] , \memory[25][53] , \memory[25][52] ,
         \memory[25][51] , \memory[25][50] , \memory[25][49] ,
         \memory[25][48] , \memory[25][47] , \memory[25][46] ,
         \memory[25][45] , \memory[25][44] , \memory[25][43] ,
         \memory[25][42] , \memory[25][41] , \memory[25][40] ,
         \memory[25][39] , \memory[25][38] , \memory[25][37] ,
         \memory[25][36] , \memory[25][35] , \memory[25][34] ,
         \memory[25][33] , \memory[25][32] , \memory[25][31] ,
         \memory[25][30] , \memory[25][29] , \memory[25][28] ,
         \memory[25][27] , \memory[25][26] , \memory[25][25] ,
         \memory[25][24] , \memory[25][23] , \memory[25][22] ,
         \memory[25][21] , \memory[25][20] , \memory[25][19] ,
         \memory[25][18] , \memory[25][17] , \memory[25][16] ,
         \memory[25][15] , \memory[25][14] , \memory[25][13] ,
         \memory[25][12] , \memory[25][11] , \memory[25][10] , \memory[25][9] ,
         \memory[25][8] , \memory[25][7] , \memory[25][6] , \memory[25][5] ,
         \memory[25][4] , \memory[25][3] , \memory[25][2] , \memory[25][1] ,
         \memory[25][0] , \memory[24][70] , \memory[24][69] , \memory[24][68] ,
         \memory[24][67] , \memory[24][66] , \memory[24][65] ,
         \memory[24][64] , \memory[24][63] , \memory[24][62] ,
         \memory[24][61] , \memory[24][60] , \memory[24][59] ,
         \memory[24][58] , \memory[24][57] , \memory[24][56] ,
         \memory[24][55] , \memory[24][54] , \memory[24][53] ,
         \memory[24][52] , \memory[24][51] , \memory[24][50] ,
         \memory[24][49] , \memory[24][48] , \memory[24][47] ,
         \memory[24][46] , \memory[24][45] , \memory[24][44] ,
         \memory[24][43] , \memory[24][42] , \memory[24][41] ,
         \memory[24][40] , \memory[24][39] , \memory[24][38] ,
         \memory[24][37] , \memory[24][36] , \memory[24][35] ,
         \memory[24][34] , \memory[24][33] , \memory[24][32] ,
         \memory[24][31] , \memory[24][30] , \memory[24][29] ,
         \memory[24][28] , \memory[24][27] , \memory[24][26] ,
         \memory[24][25] , \memory[24][24] , \memory[24][23] ,
         \memory[24][22] , \memory[24][21] , \memory[24][20] ,
         \memory[24][19] , \memory[24][18] , \memory[24][17] ,
         \memory[24][16] , \memory[24][15] , \memory[24][14] ,
         \memory[24][13] , \memory[24][12] , \memory[24][11] ,
         \memory[24][10] , \memory[24][9] , \memory[24][8] , \memory[24][7] ,
         \memory[24][6] , \memory[24][5] , \memory[24][4] , \memory[24][3] ,
         \memory[24][2] , \memory[24][1] , \memory[24][0] , \memory[23][70] ,
         \memory[23][69] , \memory[23][68] , \memory[23][67] ,
         \memory[23][66] , \memory[23][65] , \memory[23][64] ,
         \memory[23][63] , \memory[23][62] , \memory[23][61] ,
         \memory[23][60] , \memory[23][59] , \memory[23][58] ,
         \memory[23][57] , \memory[23][56] , \memory[23][55] ,
         \memory[23][54] , \memory[23][53] , \memory[23][52] ,
         \memory[23][51] , \memory[23][50] , \memory[23][49] ,
         \memory[23][48] , \memory[23][47] , \memory[23][46] ,
         \memory[23][45] , \memory[23][44] , \memory[23][43] ,
         \memory[23][42] , \memory[23][41] , \memory[23][40] ,
         \memory[23][39] , \memory[23][38] , \memory[23][37] ,
         \memory[23][36] , \memory[23][35] , \memory[23][34] ,
         \memory[23][33] , \memory[23][32] , \memory[23][31] ,
         \memory[23][30] , \memory[23][29] , \memory[23][28] ,
         \memory[23][27] , \memory[23][26] , \memory[23][25] ,
         \memory[23][24] , \memory[23][23] , \memory[23][22] ,
         \memory[23][21] , \memory[23][20] , \memory[23][19] ,
         \memory[23][18] , \memory[23][17] , \memory[23][16] ,
         \memory[23][15] , \memory[23][14] , \memory[23][13] ,
         \memory[23][12] , \memory[23][11] , \memory[23][10] , \memory[23][9] ,
         \memory[23][8] , \memory[23][7] , \memory[23][6] , \memory[23][5] ,
         \memory[23][4] , \memory[23][3] , \memory[23][2] , \memory[23][1] ,
         \memory[23][0] , \memory[22][70] , \memory[22][69] , \memory[22][68] ,
         \memory[22][67] , \memory[22][66] , \memory[22][65] ,
         \memory[22][64] , \memory[22][63] , \memory[22][62] ,
         \memory[22][61] , \memory[22][60] , \memory[22][59] ,
         \memory[22][58] , \memory[22][57] , \memory[22][56] ,
         \memory[22][55] , \memory[22][54] , \memory[22][53] ,
         \memory[22][52] , \memory[22][51] , \memory[22][50] ,
         \memory[22][49] , \memory[22][48] , \memory[22][47] ,
         \memory[22][46] , \memory[22][45] , \memory[22][44] ,
         \memory[22][43] , \memory[22][42] , \memory[22][41] ,
         \memory[22][40] , \memory[22][39] , \memory[22][38] ,
         \memory[22][37] , \memory[22][36] , \memory[22][35] ,
         \memory[22][34] , \memory[22][33] , \memory[22][32] ,
         \memory[22][31] , \memory[22][30] , \memory[22][29] ,
         \memory[22][28] , \memory[22][27] , \memory[22][26] ,
         \memory[22][25] , \memory[22][24] , \memory[22][23] ,
         \memory[22][22] , \memory[22][21] , \memory[22][20] ,
         \memory[22][19] , \memory[22][18] , \memory[22][17] ,
         \memory[22][16] , \memory[22][15] , \memory[22][14] ,
         \memory[22][13] , \memory[22][12] , \memory[22][11] ,
         \memory[22][10] , \memory[22][9] , \memory[22][8] , \memory[22][7] ,
         \memory[22][6] , \memory[22][5] , \memory[22][4] , \memory[22][3] ,
         \memory[22][2] , \memory[22][1] , \memory[22][0] , \memory[21][70] ,
         \memory[21][69] , \memory[21][68] , \memory[21][67] ,
         \memory[21][66] , \memory[21][65] , \memory[21][64] ,
         \memory[21][63] , \memory[21][62] , \memory[21][61] ,
         \memory[21][60] , \memory[21][59] , \memory[21][58] ,
         \memory[21][57] , \memory[21][56] , \memory[21][55] ,
         \memory[21][54] , \memory[21][53] , \memory[21][52] ,
         \memory[21][51] , \memory[21][50] , \memory[21][49] ,
         \memory[21][48] , \memory[21][47] , \memory[21][46] ,
         \memory[21][45] , \memory[21][44] , \memory[21][43] ,
         \memory[21][42] , \memory[21][41] , \memory[21][40] ,
         \memory[21][39] , \memory[21][38] , \memory[21][37] ,
         \memory[21][36] , \memory[21][35] , \memory[21][34] ,
         \memory[21][33] , \memory[21][32] , \memory[21][31] ,
         \memory[21][30] , \memory[21][29] , \memory[21][28] ,
         \memory[21][27] , \memory[21][26] , \memory[21][25] ,
         \memory[21][24] , \memory[21][23] , \memory[21][22] ,
         \memory[21][21] , \memory[21][20] , \memory[21][19] ,
         \memory[21][18] , \memory[21][17] , \memory[21][16] ,
         \memory[21][15] , \memory[21][14] , \memory[21][13] ,
         \memory[21][12] , \memory[21][11] , \memory[21][10] , \memory[21][9] ,
         \memory[21][8] , \memory[21][7] , \memory[21][6] , \memory[21][5] ,
         \memory[21][4] , \memory[21][3] , \memory[21][2] , \memory[21][1] ,
         \memory[21][0] , \memory[20][70] , \memory[20][69] , \memory[20][68] ,
         \memory[20][67] , \memory[20][66] , \memory[20][65] ,
         \memory[20][64] , \memory[20][63] , \memory[20][62] ,
         \memory[20][61] , \memory[20][60] , \memory[20][59] ,
         \memory[20][58] , \memory[20][57] , \memory[20][56] ,
         \memory[20][55] , \memory[20][54] , \memory[20][53] ,
         \memory[20][52] , \memory[20][51] , \memory[20][50] ,
         \memory[20][49] , \memory[20][48] , \memory[20][47] ,
         \memory[20][46] , \memory[20][45] , \memory[20][44] ,
         \memory[20][43] , \memory[20][42] , \memory[20][41] ,
         \memory[20][40] , \memory[20][39] , \memory[20][38] ,
         \memory[20][37] , \memory[20][36] , \memory[20][35] ,
         \memory[20][34] , \memory[20][33] , \memory[20][32] ,
         \memory[20][31] , \memory[20][30] , \memory[20][29] ,
         \memory[20][28] , \memory[20][27] , \memory[20][26] ,
         \memory[20][25] , \memory[20][24] , \memory[20][23] ,
         \memory[20][22] , \memory[20][21] , \memory[20][20] ,
         \memory[20][19] , \memory[20][18] , \memory[20][17] ,
         \memory[20][16] , \memory[20][15] , \memory[20][14] ,
         \memory[20][13] , \memory[20][12] , \memory[20][11] ,
         \memory[20][10] , \memory[20][9] , \memory[20][8] , \memory[20][7] ,
         \memory[20][6] , \memory[20][5] , \memory[20][4] , \memory[20][3] ,
         \memory[20][2] , \memory[20][1] , \memory[20][0] , \memory[19][70] ,
         \memory[19][69] , \memory[19][68] , \memory[19][67] ,
         \memory[19][66] , \memory[19][65] , \memory[19][64] ,
         \memory[19][63] , \memory[19][62] , \memory[19][61] ,
         \memory[19][60] , \memory[19][59] , \memory[19][58] ,
         \memory[19][57] , \memory[19][56] , \memory[19][55] ,
         \memory[19][54] , \memory[19][53] , \memory[19][52] ,
         \memory[19][51] , \memory[19][50] , \memory[19][49] ,
         \memory[19][48] , \memory[19][47] , \memory[19][46] ,
         \memory[19][45] , \memory[19][44] , \memory[19][43] ,
         \memory[19][42] , \memory[19][41] , \memory[19][40] ,
         \memory[19][39] , \memory[19][38] , \memory[19][37] ,
         \memory[19][36] , \memory[19][35] , \memory[19][34] ,
         \memory[19][33] , \memory[19][32] , \memory[19][31] ,
         \memory[19][30] , \memory[19][29] , \memory[19][28] ,
         \memory[19][27] , \memory[19][26] , \memory[19][25] ,
         \memory[19][24] , \memory[19][23] , \memory[19][22] ,
         \memory[19][21] , \memory[19][20] , \memory[19][19] ,
         \memory[19][18] , \memory[19][17] , \memory[19][16] ,
         \memory[19][15] , \memory[19][14] , \memory[19][13] ,
         \memory[19][12] , \memory[19][11] , \memory[19][10] , \memory[19][9] ,
         \memory[19][8] , \memory[19][7] , \memory[19][6] , \memory[19][5] ,
         \memory[19][4] , \memory[19][3] , \memory[19][2] , \memory[19][1] ,
         \memory[19][0] , \memory[18][70] , \memory[18][69] , \memory[18][68] ,
         \memory[18][67] , \memory[18][66] , \memory[18][65] ,
         \memory[18][64] , \memory[18][63] , \memory[18][62] ,
         \memory[18][61] , \memory[18][60] , \memory[18][59] ,
         \memory[18][58] , \memory[18][57] , \memory[18][56] ,
         \memory[18][55] , \memory[18][54] , \memory[18][53] ,
         \memory[18][52] , \memory[18][51] , \memory[18][50] ,
         \memory[18][49] , \memory[18][48] , \memory[18][47] ,
         \memory[18][46] , \memory[18][45] , \memory[18][44] ,
         \memory[18][43] , \memory[18][42] , \memory[18][41] ,
         \memory[18][40] , \memory[18][39] , \memory[18][38] ,
         \memory[18][37] , \memory[18][36] , \memory[18][35] ,
         \memory[18][34] , \memory[18][33] , \memory[18][32] ,
         \memory[18][31] , \memory[18][30] , \memory[18][29] ,
         \memory[18][28] , \memory[18][27] , \memory[18][26] ,
         \memory[18][25] , \memory[18][24] , \memory[18][23] ,
         \memory[18][22] , \memory[18][21] , \memory[18][20] ,
         \memory[18][19] , \memory[18][18] , \memory[18][17] ,
         \memory[18][16] , \memory[18][15] , \memory[18][14] ,
         \memory[18][13] , \memory[18][12] , \memory[18][11] ,
         \memory[18][10] , \memory[18][9] , \memory[18][8] , \memory[18][7] ,
         \memory[18][6] , \memory[18][5] , \memory[18][4] , \memory[18][3] ,
         \memory[18][2] , \memory[18][1] , \memory[18][0] , \memory[17][70] ,
         \memory[17][69] , \memory[17][68] , \memory[17][67] ,
         \memory[17][66] , \memory[17][65] , \memory[17][64] ,
         \memory[17][63] , \memory[17][62] , \memory[17][61] ,
         \memory[17][60] , \memory[17][59] , \memory[17][58] ,
         \memory[17][57] , \memory[17][56] , \memory[17][55] ,
         \memory[17][54] , \memory[17][53] , \memory[17][52] ,
         \memory[17][51] , \memory[17][50] , \memory[17][49] ,
         \memory[17][48] , \memory[17][47] , \memory[17][46] ,
         \memory[17][45] , \memory[17][44] , \memory[17][43] ,
         \memory[17][42] , \memory[17][41] , \memory[17][40] ,
         \memory[17][39] , \memory[17][38] , \memory[17][37] ,
         \memory[17][36] , \memory[17][35] , \memory[17][34] ,
         \memory[17][33] , \memory[17][32] , \memory[17][31] ,
         \memory[17][30] , \memory[17][29] , \memory[17][28] ,
         \memory[17][27] , \memory[17][26] , \memory[17][25] ,
         \memory[17][24] , \memory[17][23] , \memory[17][22] ,
         \memory[17][21] , \memory[17][20] , \memory[17][19] ,
         \memory[17][18] , \memory[17][17] , \memory[17][16] ,
         \memory[17][15] , \memory[17][14] , \memory[17][13] ,
         \memory[17][12] , \memory[17][11] , \memory[17][10] , \memory[17][9] ,
         \memory[17][8] , \memory[17][7] , \memory[17][6] , \memory[17][5] ,
         \memory[17][4] , \memory[17][3] , \memory[17][2] , \memory[17][1] ,
         \memory[17][0] , \memory[16][70] , \memory[16][69] , \memory[16][68] ,
         \memory[16][67] , \memory[16][66] , \memory[16][65] ,
         \memory[16][64] , \memory[16][63] , \memory[16][62] ,
         \memory[16][61] , \memory[16][60] , \memory[16][59] ,
         \memory[16][58] , \memory[16][57] , \memory[16][56] ,
         \memory[16][55] , \memory[16][54] , \memory[16][53] ,
         \memory[16][52] , \memory[16][51] , \memory[16][50] ,
         \memory[16][49] , \memory[16][48] , \memory[16][47] ,
         \memory[16][46] , \memory[16][45] , \memory[16][44] ,
         \memory[16][43] , \memory[16][42] , \memory[16][41] ,
         \memory[16][40] , \memory[16][39] , \memory[16][38] ,
         \memory[16][37] , \memory[16][36] , \memory[16][35] ,
         \memory[16][34] , \memory[16][33] , \memory[16][32] ,
         \memory[16][31] , \memory[16][30] , \memory[16][29] ,
         \memory[16][28] , \memory[16][27] , \memory[16][26] ,
         \memory[16][25] , \memory[16][24] , \memory[16][23] ,
         \memory[16][22] , \memory[16][21] , \memory[16][20] ,
         \memory[16][19] , \memory[16][18] , \memory[16][17] ,
         \memory[16][16] , \memory[16][15] , \memory[16][14] ,
         \memory[16][13] , \memory[16][12] , \memory[16][11] ,
         \memory[16][10] , \memory[16][9] , \memory[16][8] , \memory[16][7] ,
         \memory[16][6] , \memory[16][5] , \memory[16][4] , \memory[16][3] ,
         \memory[16][2] , \memory[16][1] , \memory[16][0] , \memory[15][70] ,
         \memory[15][69] , \memory[15][68] , \memory[15][67] ,
         \memory[15][66] , \memory[15][65] , \memory[15][64] ,
         \memory[15][63] , \memory[15][62] , \memory[15][61] ,
         \memory[15][60] , \memory[15][59] , \memory[15][58] ,
         \memory[15][57] , \memory[15][56] , \memory[15][55] ,
         \memory[15][54] , \memory[15][53] , \memory[15][52] ,
         \memory[15][51] , \memory[15][50] , \memory[15][49] ,
         \memory[15][48] , \memory[15][47] , \memory[15][46] ,
         \memory[15][45] , \memory[15][44] , \memory[15][43] ,
         \memory[15][42] , \memory[15][41] , \memory[15][40] ,
         \memory[15][39] , \memory[15][38] , \memory[15][37] ,
         \memory[15][36] , \memory[15][35] , \memory[15][34] ,
         \memory[15][33] , \memory[15][32] , \memory[15][31] ,
         \memory[15][30] , \memory[15][29] , \memory[15][28] ,
         \memory[15][27] , \memory[15][26] , \memory[15][25] ,
         \memory[15][24] , \memory[15][23] , \memory[15][22] ,
         \memory[15][21] , \memory[15][20] , \memory[15][19] ,
         \memory[15][18] , \memory[15][17] , \memory[15][16] ,
         \memory[15][15] , \memory[15][14] , \memory[15][13] ,
         \memory[15][12] , \memory[15][11] , \memory[15][10] , \memory[15][9] ,
         \memory[15][8] , \memory[15][7] , \memory[15][6] , \memory[15][5] ,
         \memory[15][4] , \memory[15][3] , \memory[15][2] , \memory[15][1] ,
         \memory[15][0] , \memory[14][70] , \memory[14][69] , \memory[14][68] ,
         \memory[14][67] , \memory[14][66] , \memory[14][65] ,
         \memory[14][64] , \memory[14][63] , \memory[14][62] ,
         \memory[14][61] , \memory[14][60] , \memory[14][59] ,
         \memory[14][58] , \memory[14][57] , \memory[14][56] ,
         \memory[14][55] , \memory[14][54] , \memory[14][53] ,
         \memory[14][52] , \memory[14][51] , \memory[14][50] ,
         \memory[14][49] , \memory[14][48] , \memory[14][47] ,
         \memory[14][46] , \memory[14][45] , \memory[14][44] ,
         \memory[14][43] , \memory[14][42] , \memory[14][41] ,
         \memory[14][40] , \memory[14][39] , \memory[14][38] ,
         \memory[14][37] , \memory[14][36] , \memory[14][35] ,
         \memory[14][34] , \memory[14][33] , \memory[14][32] ,
         \memory[14][31] , \memory[14][30] , \memory[14][29] ,
         \memory[14][28] , \memory[14][27] , \memory[14][26] ,
         \memory[14][25] , \memory[14][24] , \memory[14][23] ,
         \memory[14][22] , \memory[14][21] , \memory[14][20] ,
         \memory[14][19] , \memory[14][18] , \memory[14][17] ,
         \memory[14][16] , \memory[14][15] , \memory[14][14] ,
         \memory[14][13] , \memory[14][12] , \memory[14][11] ,
         \memory[14][10] , \memory[14][9] , \memory[14][8] , \memory[14][7] ,
         \memory[14][6] , \memory[14][5] , \memory[14][4] , \memory[14][3] ,
         \memory[14][2] , \memory[14][1] , \memory[14][0] , \memory[13][70] ,
         \memory[13][69] , \memory[13][68] , \memory[13][67] ,
         \memory[13][66] , \memory[13][65] , \memory[13][64] ,
         \memory[13][63] , \memory[13][62] , \memory[13][61] ,
         \memory[13][60] , \memory[13][59] , \memory[13][58] ,
         \memory[13][57] , \memory[13][56] , \memory[13][55] ,
         \memory[13][54] , \memory[13][53] , \memory[13][52] ,
         \memory[13][51] , \memory[13][50] , \memory[13][49] ,
         \memory[13][48] , \memory[13][47] , \memory[13][46] ,
         \memory[13][45] , \memory[13][44] , \memory[13][43] ,
         \memory[13][42] , \memory[13][41] , \memory[13][40] ,
         \memory[13][39] , \memory[13][38] , \memory[13][37] ,
         \memory[13][36] , \memory[13][35] , \memory[13][34] ,
         \memory[13][33] , \memory[13][32] , \memory[13][31] ,
         \memory[13][30] , \memory[13][29] , \memory[13][28] ,
         \memory[13][27] , \memory[13][26] , \memory[13][25] ,
         \memory[13][24] , \memory[13][23] , \memory[13][22] ,
         \memory[13][21] , \memory[13][20] , \memory[13][19] ,
         \memory[13][18] , \memory[13][17] , \memory[13][16] ,
         \memory[13][15] , \memory[13][14] , \memory[13][13] ,
         \memory[13][12] , \memory[13][11] , \memory[13][10] , \memory[13][9] ,
         \memory[13][8] , \memory[13][7] , \memory[13][6] , \memory[13][5] ,
         \memory[13][4] , \memory[13][3] , \memory[13][2] , \memory[13][1] ,
         \memory[13][0] , \memory[12][70] , \memory[12][69] , \memory[12][68] ,
         \memory[12][67] , \memory[12][66] , \memory[12][65] ,
         \memory[12][64] , \memory[12][63] , \memory[12][62] ,
         \memory[12][61] , \memory[12][60] , \memory[12][59] ,
         \memory[12][58] , \memory[12][57] , \memory[12][56] ,
         \memory[12][55] , \memory[12][54] , \memory[12][53] ,
         \memory[12][52] , \memory[12][51] , \memory[12][50] ,
         \memory[12][49] , \memory[12][48] , \memory[12][47] ,
         \memory[12][46] , \memory[12][45] , \memory[12][44] ,
         \memory[12][43] , \memory[12][42] , \memory[12][41] ,
         \memory[12][40] , \memory[12][39] , \memory[12][38] ,
         \memory[12][37] , \memory[12][36] , \memory[12][35] ,
         \memory[12][34] , \memory[12][33] , \memory[12][32] ,
         \memory[12][31] , \memory[12][30] , \memory[12][29] ,
         \memory[12][28] , \memory[12][27] , \memory[12][26] ,
         \memory[12][25] , \memory[12][24] , \memory[12][23] ,
         \memory[12][22] , \memory[12][21] , \memory[12][20] ,
         \memory[12][19] , \memory[12][18] , \memory[12][17] ,
         \memory[12][16] , \memory[12][15] , \memory[12][14] ,
         \memory[12][13] , \memory[12][12] , \memory[12][11] ,
         \memory[12][10] , \memory[12][9] , \memory[12][8] , \memory[12][7] ,
         \memory[12][6] , \memory[12][5] , \memory[12][4] , \memory[12][3] ,
         \memory[12][2] , \memory[12][1] , \memory[12][0] , \memory[11][70] ,
         \memory[11][69] , \memory[11][68] , \memory[11][67] ,
         \memory[11][66] , \memory[11][65] , \memory[11][64] ,
         \memory[11][63] , \memory[11][62] , \memory[11][61] ,
         \memory[11][60] , \memory[11][59] , \memory[11][58] ,
         \memory[11][57] , \memory[11][56] , \memory[11][55] ,
         \memory[11][54] , \memory[11][53] , \memory[11][52] ,
         \memory[11][51] , \memory[11][50] , \memory[11][49] ,
         \memory[11][48] , \memory[11][47] , \memory[11][46] ,
         \memory[11][45] , \memory[11][44] , \memory[11][43] ,
         \memory[11][42] , \memory[11][41] , \memory[11][40] ,
         \memory[11][39] , \memory[11][38] , \memory[11][37] ,
         \memory[11][36] , \memory[11][35] , \memory[11][34] ,
         \memory[11][33] , \memory[11][32] , \memory[11][31] ,
         \memory[11][30] , \memory[11][29] , \memory[11][28] ,
         \memory[11][27] , \memory[11][26] , \memory[11][25] ,
         \memory[11][24] , \memory[11][23] , \memory[11][22] ,
         \memory[11][21] , \memory[11][20] , \memory[11][19] ,
         \memory[11][18] , \memory[11][17] , \memory[11][16] ,
         \memory[11][15] , \memory[11][14] , \memory[11][13] ,
         \memory[11][12] , \memory[11][11] , \memory[11][10] , \memory[11][9] ,
         \memory[11][8] , \memory[11][7] , \memory[11][6] , \memory[11][5] ,
         \memory[11][4] , \memory[11][3] , \memory[11][2] , \memory[11][1] ,
         \memory[11][0] , \memory[10][70] , \memory[10][69] , \memory[10][68] ,
         \memory[10][67] , \memory[10][66] , \memory[10][65] ,
         \memory[10][64] , \memory[10][63] , \memory[10][62] ,
         \memory[10][61] , \memory[10][60] , \memory[10][59] ,
         \memory[10][58] , \memory[10][57] , \memory[10][56] ,
         \memory[10][55] , \memory[10][54] , \memory[10][53] ,
         \memory[10][52] , \memory[10][51] , \memory[10][50] ,
         \memory[10][49] , \memory[10][48] , \memory[10][47] ,
         \memory[10][46] , \memory[10][45] , \memory[10][44] ,
         \memory[10][43] , \memory[10][42] , \memory[10][41] ,
         \memory[10][40] , \memory[10][39] , \memory[10][38] ,
         \memory[10][37] , \memory[10][36] , \memory[10][35] ,
         \memory[10][34] , \memory[10][33] , \memory[10][32] ,
         \memory[10][31] , \memory[10][30] , \memory[10][29] ,
         \memory[10][28] , \memory[10][27] , \memory[10][26] ,
         \memory[10][25] , \memory[10][24] , \memory[10][23] ,
         \memory[10][22] , \memory[10][21] , \memory[10][20] ,
         \memory[10][19] , \memory[10][18] , \memory[10][17] ,
         \memory[10][16] , \memory[10][15] , \memory[10][14] ,
         \memory[10][13] , \memory[10][12] , \memory[10][11] ,
         \memory[10][10] , \memory[10][9] , \memory[10][8] , \memory[10][7] ,
         \memory[10][6] , \memory[10][5] , \memory[10][4] , \memory[10][3] ,
         \memory[10][2] , \memory[10][1] , \memory[10][0] , \memory[9][70] ,
         \memory[9][69] , \memory[9][68] , \memory[9][67] , \memory[9][66] ,
         \memory[9][65] , \memory[9][64] , \memory[9][63] , \memory[9][62] ,
         \memory[9][61] , \memory[9][60] , \memory[9][59] , \memory[9][58] ,
         \memory[9][57] , \memory[9][56] , \memory[9][55] , \memory[9][54] ,
         \memory[9][53] , \memory[9][52] , \memory[9][51] , \memory[9][50] ,
         \memory[9][49] , \memory[9][48] , \memory[9][47] , \memory[9][46] ,
         \memory[9][45] , \memory[9][44] , \memory[9][43] , \memory[9][42] ,
         \memory[9][41] , \memory[9][40] , \memory[9][39] , \memory[9][38] ,
         \memory[9][37] , \memory[9][36] , \memory[9][35] , \memory[9][34] ,
         \memory[9][33] , \memory[9][32] , \memory[9][31] , \memory[9][30] ,
         \memory[9][29] , \memory[9][28] , \memory[9][27] , \memory[9][26] ,
         \memory[9][25] , \memory[9][24] , \memory[9][23] , \memory[9][22] ,
         \memory[9][21] , \memory[9][20] , \memory[9][19] , \memory[9][18] ,
         \memory[9][17] , \memory[9][16] , \memory[9][15] , \memory[9][14] ,
         \memory[9][13] , \memory[9][12] , \memory[9][11] , \memory[9][10] ,
         \memory[9][9] , \memory[9][8] , \memory[9][7] , \memory[9][6] ,
         \memory[9][5] , \memory[9][4] , \memory[9][3] , \memory[9][2] ,
         \memory[9][1] , \memory[9][0] , \memory[8][70] , \memory[8][69] ,
         \memory[8][68] , \memory[8][67] , \memory[8][66] , \memory[8][65] ,
         \memory[8][64] , \memory[8][63] , \memory[8][62] , \memory[8][61] ,
         \memory[8][60] , \memory[8][59] , \memory[8][58] , \memory[8][57] ,
         \memory[8][56] , \memory[8][55] , \memory[8][54] , \memory[8][53] ,
         \memory[8][52] , \memory[8][51] , \memory[8][50] , \memory[8][49] ,
         \memory[8][48] , \memory[8][47] , \memory[8][46] , \memory[8][45] ,
         \memory[8][44] , \memory[8][43] , \memory[8][42] , \memory[8][41] ,
         \memory[8][40] , \memory[8][39] , \memory[8][38] , \memory[8][37] ,
         \memory[8][36] , \memory[8][35] , \memory[8][34] , \memory[8][33] ,
         \memory[8][32] , \memory[8][31] , \memory[8][30] , \memory[8][29] ,
         \memory[8][28] , \memory[8][27] , \memory[8][26] , \memory[8][25] ,
         \memory[8][24] , \memory[8][23] , \memory[8][22] , \memory[8][21] ,
         \memory[8][20] , \memory[8][19] , \memory[8][18] , \memory[8][17] ,
         \memory[8][16] , \memory[8][15] , \memory[8][14] , \memory[8][13] ,
         \memory[8][12] , \memory[8][11] , \memory[8][10] , \memory[8][9] ,
         \memory[8][8] , \memory[8][7] , \memory[8][6] , \memory[8][5] ,
         \memory[8][4] , \memory[8][3] , \memory[8][2] , \memory[8][1] ,
         \memory[8][0] , \memory[7][70] , \memory[7][69] , \memory[7][68] ,
         \memory[7][67] , \memory[7][66] , \memory[7][65] , \memory[7][64] ,
         \memory[7][63] , \memory[7][62] , \memory[7][61] , \memory[7][60] ,
         \memory[7][59] , \memory[7][58] , \memory[7][57] , \memory[7][56] ,
         \memory[7][55] , \memory[7][54] , \memory[7][53] , \memory[7][52] ,
         \memory[7][51] , \memory[7][50] , \memory[7][49] , \memory[7][48] ,
         \memory[7][47] , \memory[7][46] , \memory[7][45] , \memory[7][44] ,
         \memory[7][43] , \memory[7][42] , \memory[7][41] , \memory[7][40] ,
         \memory[7][39] , \memory[7][38] , \memory[7][37] , \memory[7][36] ,
         \memory[7][35] , \memory[7][34] , \memory[7][33] , \memory[7][32] ,
         \memory[7][31] , \memory[7][30] , \memory[7][29] , \memory[7][28] ,
         \memory[7][27] , \memory[7][26] , \memory[7][25] , \memory[7][24] ,
         \memory[7][23] , \memory[7][22] , \memory[7][21] , \memory[7][20] ,
         \memory[7][19] , \memory[7][18] , \memory[7][17] , \memory[7][16] ,
         \memory[7][15] , \memory[7][14] , \memory[7][13] , \memory[7][12] ,
         \memory[7][11] , \memory[7][10] , \memory[7][9] , \memory[7][8] ,
         \memory[7][7] , \memory[7][6] , \memory[7][5] , \memory[7][4] ,
         \memory[7][3] , \memory[7][2] , \memory[7][1] , \memory[7][0] ,
         \memory[6][70] , \memory[6][69] , \memory[6][68] , \memory[6][67] ,
         \memory[6][66] , \memory[6][65] , \memory[6][64] , \memory[6][63] ,
         \memory[6][62] , \memory[6][61] , \memory[6][60] , \memory[6][59] ,
         \memory[6][58] , \memory[6][57] , \memory[6][56] , \memory[6][55] ,
         \memory[6][54] , \memory[6][53] , \memory[6][52] , \memory[6][51] ,
         \memory[6][50] , \memory[6][49] , \memory[6][48] , \memory[6][47] ,
         \memory[6][46] , \memory[6][45] , \memory[6][44] , \memory[6][43] ,
         \memory[6][42] , \memory[6][41] , \memory[6][40] , \memory[6][39] ,
         \memory[6][38] , \memory[6][37] , \memory[6][36] , \memory[6][35] ,
         \memory[6][34] , \memory[6][33] , \memory[6][32] , \memory[6][31] ,
         \memory[6][30] , \memory[6][29] , \memory[6][28] , \memory[6][27] ,
         \memory[6][26] , \memory[6][25] , \memory[6][24] , \memory[6][23] ,
         \memory[6][22] , \memory[6][21] , \memory[6][20] , \memory[6][19] ,
         \memory[6][18] , \memory[6][17] , \memory[6][16] , \memory[6][15] ,
         \memory[6][14] , \memory[6][13] , \memory[6][12] , \memory[6][11] ,
         \memory[6][10] , \memory[6][9] , \memory[6][8] , \memory[6][7] ,
         \memory[6][6] , \memory[6][5] , \memory[6][4] , \memory[6][3] ,
         \memory[6][2] , \memory[6][1] , \memory[6][0] , \memory[5][70] ,
         \memory[5][69] , \memory[5][68] , \memory[5][67] , \memory[5][66] ,
         \memory[5][65] , \memory[5][64] , \memory[5][63] , \memory[5][62] ,
         \memory[5][61] , \memory[5][60] , \memory[5][59] , \memory[5][58] ,
         \memory[5][57] , \memory[5][56] , \memory[5][55] , \memory[5][54] ,
         \memory[5][53] , \memory[5][52] , \memory[5][51] , \memory[5][50] ,
         \memory[5][49] , \memory[5][48] , \memory[5][47] , \memory[5][46] ,
         \memory[5][45] , \memory[5][44] , \memory[5][43] , \memory[5][42] ,
         \memory[5][41] , \memory[5][40] , \memory[5][39] , \memory[5][38] ,
         \memory[5][37] , \memory[5][36] , \memory[5][35] , \memory[5][34] ,
         \memory[5][33] , \memory[5][32] , \memory[5][31] , \memory[5][30] ,
         \memory[5][29] , \memory[5][28] , \memory[5][27] , \memory[5][26] ,
         \memory[5][25] , \memory[5][24] , \memory[5][23] , \memory[5][22] ,
         \memory[5][21] , \memory[5][20] , \memory[5][19] , \memory[5][18] ,
         \memory[5][17] , \memory[5][16] , \memory[5][15] , \memory[5][14] ,
         \memory[5][13] , \memory[5][12] , \memory[5][11] , \memory[5][10] ,
         \memory[5][9] , \memory[5][8] , \memory[5][7] , \memory[5][6] ,
         \memory[5][5] , \memory[5][4] , \memory[5][3] , \memory[5][2] ,
         \memory[5][1] , \memory[5][0] , \memory[4][70] , \memory[4][69] ,
         \memory[4][68] , \memory[4][67] , \memory[4][66] , \memory[4][65] ,
         \memory[4][64] , \memory[4][63] , \memory[4][62] , \memory[4][61] ,
         \memory[4][60] , \memory[4][59] , \memory[4][58] , \memory[4][57] ,
         \memory[4][56] , \memory[4][55] , \memory[4][54] , \memory[4][53] ,
         \memory[4][52] , \memory[4][51] , \memory[4][50] , \memory[4][49] ,
         \memory[4][48] , \memory[4][47] , \memory[4][46] , \memory[4][45] ,
         \memory[4][44] , \memory[4][43] , \memory[4][42] , \memory[4][41] ,
         \memory[4][40] , \memory[4][39] , \memory[4][38] , \memory[4][37] ,
         \memory[4][36] , \memory[4][35] , \memory[4][34] , \memory[4][33] ,
         \memory[4][32] , \memory[4][31] , \memory[4][30] , \memory[4][29] ,
         \memory[4][28] , \memory[4][27] , \memory[4][26] , \memory[4][25] ,
         \memory[4][24] , \memory[4][23] , \memory[4][22] , \memory[4][21] ,
         \memory[4][20] , \memory[4][19] , \memory[4][18] , \memory[4][17] ,
         \memory[4][16] , \memory[4][15] , \memory[4][14] , \memory[4][13] ,
         \memory[4][12] , \memory[4][11] , \memory[4][10] , \memory[4][9] ,
         \memory[4][8] , \memory[4][7] , \memory[4][6] , \memory[4][5] ,
         \memory[4][4] , \memory[4][3] , \memory[4][2] , \memory[4][1] ,
         \memory[4][0] , \memory[3][70] , \memory[3][69] , \memory[3][68] ,
         \memory[3][67] , \memory[3][66] , \memory[3][65] , \memory[3][64] ,
         \memory[3][63] , \memory[3][62] , \memory[3][61] , \memory[3][60] ,
         \memory[3][59] , \memory[3][58] , \memory[3][57] , \memory[3][56] ,
         \memory[3][55] , \memory[3][54] , \memory[3][53] , \memory[3][52] ,
         \memory[3][51] , \memory[3][50] , \memory[3][49] , \memory[3][48] ,
         \memory[3][47] , \memory[3][46] , \memory[3][45] , \memory[3][44] ,
         \memory[3][43] , \memory[3][42] , \memory[3][41] , \memory[3][40] ,
         \memory[3][39] , \memory[3][38] , \memory[3][37] , \memory[3][36] ,
         \memory[3][35] , \memory[3][34] , \memory[3][33] , \memory[3][32] ,
         \memory[3][31] , \memory[3][30] , \memory[3][29] , \memory[3][28] ,
         \memory[3][27] , \memory[3][26] , \memory[3][25] , \memory[3][24] ,
         \memory[3][23] , \memory[3][22] , \memory[3][21] , \memory[3][20] ,
         \memory[3][19] , \memory[3][18] , \memory[3][17] , \memory[3][16] ,
         \memory[3][15] , \memory[3][14] , \memory[3][13] , \memory[3][12] ,
         \memory[3][11] , \memory[3][10] , \memory[3][9] , \memory[3][8] ,
         \memory[3][7] , \memory[3][6] , \memory[3][5] , \memory[3][4] ,
         \memory[3][3] , \memory[3][2] , \memory[3][1] , \memory[3][0] ,
         \memory[2][70] , \memory[2][69] , \memory[2][68] , \memory[2][67] ,
         \memory[2][66] , \memory[2][65] , \memory[2][64] , \memory[2][63] ,
         \memory[2][62] , \memory[2][61] , \memory[2][60] , \memory[2][59] ,
         \memory[2][58] , \memory[2][57] , \memory[2][56] , \memory[2][55] ,
         \memory[2][54] , \memory[2][53] , \memory[2][52] , \memory[2][51] ,
         \memory[2][50] , \memory[2][49] , \memory[2][48] , \memory[2][47] ,
         \memory[2][46] , \memory[2][45] , \memory[2][44] , \memory[2][43] ,
         \memory[2][42] , \memory[2][41] , \memory[2][40] , \memory[2][39] ,
         \memory[2][38] , \memory[2][37] , \memory[2][36] , \memory[2][35] ,
         \memory[2][34] , \memory[2][33] , \memory[2][32] , \memory[2][31] ,
         \memory[2][30] , \memory[2][29] , \memory[2][28] , \memory[2][27] ,
         \memory[2][26] , \memory[2][25] , \memory[2][24] , \memory[2][23] ,
         \memory[2][22] , \memory[2][21] , \memory[2][20] , \memory[2][19] ,
         \memory[2][18] , \memory[2][17] , \memory[2][16] , \memory[2][15] ,
         \memory[2][14] , \memory[2][13] , \memory[2][12] , \memory[2][11] ,
         \memory[2][10] , \memory[2][9] , \memory[2][8] , \memory[2][7] ,
         \memory[2][6] , \memory[2][5] , \memory[2][4] , \memory[2][3] ,
         \memory[2][2] , \memory[2][1] , \memory[2][0] , \memory[1][70] ,
         \memory[1][69] , \memory[1][68] , \memory[1][67] , \memory[1][66] ,
         \memory[1][65] , \memory[1][64] , \memory[1][63] , \memory[1][62] ,
         \memory[1][61] , \memory[1][60] , \memory[1][59] , \memory[1][58] ,
         \memory[1][57] , \memory[1][56] , \memory[1][55] , \memory[1][54] ,
         \memory[1][53] , \memory[1][52] , \memory[1][51] , \memory[1][50] ,
         \memory[1][49] , \memory[1][48] , \memory[1][47] , \memory[1][46] ,
         \memory[1][45] , \memory[1][44] , \memory[1][43] , \memory[1][42] ,
         \memory[1][41] , \memory[1][40] , \memory[1][39] , \memory[1][38] ,
         \memory[1][37] , \memory[1][36] , \memory[1][35] , \memory[1][34] ,
         \memory[1][33] , \memory[1][32] , \memory[1][31] , \memory[1][30] ,
         \memory[1][29] , \memory[1][28] , \memory[1][27] , \memory[1][26] ,
         \memory[1][25] , \memory[1][24] , \memory[1][23] , \memory[1][22] ,
         \memory[1][21] , \memory[1][20] , \memory[1][19] , \memory[1][18] ,
         \memory[1][17] , \memory[1][16] , \memory[1][15] , \memory[1][14] ,
         \memory[1][13] , \memory[1][12] , \memory[1][11] , \memory[1][10] ,
         \memory[1][9] , \memory[1][8] , \memory[1][7] , \memory[1][6] ,
         \memory[1][5] , \memory[1][4] , \memory[1][3] , \memory[1][2] ,
         \memory[1][1] , \memory[1][0] , \memory[0][70] , \memory[0][69] ,
         \memory[0][68] , \memory[0][67] , \memory[0][66] , \memory[0][65] ,
         \memory[0][64] , \memory[0][63] , \memory[0][62] , \memory[0][61] ,
         \memory[0][60] , \memory[0][59] , \memory[0][58] , \memory[0][57] ,
         \memory[0][56] , \memory[0][55] , \memory[0][54] , \memory[0][53] ,
         \memory[0][52] , \memory[0][51] , \memory[0][50] , \memory[0][49] ,
         \memory[0][48] , \memory[0][47] , \memory[0][46] , \memory[0][45] ,
         \memory[0][44] , \memory[0][43] , \memory[0][42] , \memory[0][41] ,
         \memory[0][40] , \memory[0][39] , \memory[0][38] , \memory[0][37] ,
         \memory[0][36] , \memory[0][35] , \memory[0][34] , \memory[0][33] ,
         \memory[0][32] , \memory[0][31] , \memory[0][30] , \memory[0][29] ,
         \memory[0][28] , \memory[0][27] , \memory[0][26] , \memory[0][25] ,
         \memory[0][24] , \memory[0][23] , \memory[0][22] , \memory[0][21] ,
         \memory[0][20] , \memory[0][19] , \memory[0][18] , \memory[0][17] ,
         \memory[0][16] , \memory[0][15] , \memory[0][14] , \memory[0][13] ,
         \memory[0][12] , \memory[0][11] , \memory[0][10] , \memory[0][9] ,
         \memory[0][8] , \memory[0][7] , \memory[0][6] , \memory[0][5] ,
         \memory[0][4] , \memory[0][3] , \memory[0][2] , \memory[0][1] ,
         \memory[0][0] , N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, write, full, N114, read, empty,
         N115, N121, N122, N123, N124, N126, N127, N128, N129, N130, N131,
         N132, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N213, N214, N215, N216, N217,
         N218, N220, N221, N222, N223, N230, N231, N232, N233, N234, N235,
         N242, N243, N244, N245, N246, N247, N2521, N2522, N2523, N2524, N2525,
         N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535,
         N2536, N2537, N2538, N2539, N2610, N2617, N2681, N2688, N2752, N2759,
         N2823, N2830, N2894, N2901, N2965, N2972, N3036, N3043, N3107, N3114,
         N3178, N3185, N3249, N3256, N3320, N3327, N3391, N3398, N3462, N3469,
         N3533, N3540, N3604, N3611, N3675, N3682, N3746, N3753, N3817, N3824,
         N3888, N3895, N3959, N3966, N4030, N4037, N4101, N4108, N4172, N4179,
         N4243, N4250, N4314, N4321, N4385, N4392, N4456, N4463, N4527, N4534,
         N4598, N4605, N4669, N4676, N4740, N4747, N4811, N4818, N4960, N4961,
         N4965, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113,
         N5114, N5115, N5116, N5117, N5118, N5120, N5121, N5122, N5123, N5124,
         N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, N5134,
         N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144,
         N5145, N5146, N5147, N5148, N5149, N5150, N5151, N5152, N5153, N5154,
         N5155, N5156, N5157, N5158, N5159, N5160, N5161, N5162, N5163, N5164,
         N5165, N5166, N5167, N5168, N5169, N5170, N5171, N5172, N5173, N5174,
         N5175, N5176, N5177, N5178, N5179, N5180, N5181, N5182, N5183, N5184,
         N5185, N5186, N5187, N5188, N5189, N5190, N5191, N5192, N5193, N5194,
         N5195, N5196, N5197, N5198, N5199, N5200, N5201, N5202, N5203, N5204,
         N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212, N5213, N5214,
         N5215, N5216, N5217, N5218, N5219, N5220, N5221, N5222, N5223, N5224,
         N5225, N5226, N5227, N5228, N5229, N5230, N5231, N5232, N5233, N5234,
         N5235, N5236, N5237, N5238, N5239, N5240, N5241, N5242, N5243, N5244,
         N5245, N5246, N5247, N5248, N5249, N5250, N5251, N5252, N5253, N5254,
         N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262, N5263, N5264,
         N5265, N5266, N5267, N5268, N5269, N5270, N5271, N5272, N5273, N5274,
         N5275, N5276, N5277, N5278, N5279, N5280, N5281, N5282, N5283, N5284,
         N5285, N5286, N5287, N5288, N5289, N5290, N5291, N5292, N5293, N5294,
         N5295, N5296, N5297, N5298, N5299, N5300, N5301, N5302, N5303, N5304,
         N5305, N5306, N5307, N5308, N5309, N5310, N5311, N5312, N5313, N5314,
         n2, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, \add_116/carry[5] ,
         \add_116/carry[4] , \add_116/carry[3] , \add_116/carry[2] ,
         \r184/carry[4] , \r184/carry[3] , \r184/carry[2] , \r183/carry[4] ,
         \r183/carry[3] , \r183/carry[2] , n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939;
  wire   [6:0] lout;
  wire   [62:0] out;
  wire   [4:0] write_ptr;
  wire   [63:0] out_new;
  wire   [6:0] lout_new;
  wire   [5:0] counter;

  CNIVX4 B_13 ( .A(N5112), .Z(full) );
  CNIVX4 B_12 ( .A(N5118), .Z(empty) );
  CAN2X2 C41739 ( .A(N114), .B(N115), .Z(N210) );
  CIVX2 I_41 ( .A(N121), .Z(N122) );
  CIVX2 I_37 ( .A(empty), .Z(N5314) );
  CAN2X2 C41721 ( .A(read), .B(N5314), .Z(N115) );
  CIVX2 I_36 ( .A(full), .Z(N5313) );
  CAN2X2 C41719 ( .A(write), .B(N5313), .Z(N114) );
  CAN2X2 C41707 ( .A(N5268), .B(N5280), .Z(N5312) );
  CAN2X2 C41706 ( .A(N5268), .B(N5279), .Z(N5311) );
  CAN2X2 C41705 ( .A(N5268), .B(N5278), .Z(N5310) );
  CAN2X2 C41704 ( .A(N5268), .B(N5277), .Z(N5309) );
  CAN2X2 C41703 ( .A(N5268), .B(N5276), .Z(N5308) );
  CAN2X2 C41702 ( .A(N5268), .B(N5275), .Z(N5307) );
  CAN2X2 C41701 ( .A(N5268), .B(N5274), .Z(N5306) );
  CAN2X2 C41700 ( .A(N5268), .B(N5273), .Z(N5305) );
  CAN2X2 C41699 ( .A(N5267), .B(N5280), .Z(N5304) );
  CAN2X2 C41698 ( .A(N5267), .B(N5279), .Z(N5303) );
  CAN2X2 C41697 ( .A(N5267), .B(N5278), .Z(N5302) );
  CAN2X2 C41696 ( .A(N5267), .B(N5277), .Z(N5301) );
  CAN2X2 C41695 ( .A(N5267), .B(N5276), .Z(N5300) );
  CAN2X2 C41694 ( .A(N5267), .B(N5275), .Z(N5299) );
  CAN2X2 C41693 ( .A(N5267), .B(N5274), .Z(N5298) );
  CAN2X2 C41692 ( .A(N5267), .B(N5273), .Z(N5297) );
  CAN2X2 C41691 ( .A(N5266), .B(N5280), .Z(N5296) );
  CAN2X2 C41690 ( .A(N5266), .B(N5279), .Z(N5295) );
  CAN2X2 C41689 ( .A(N5266), .B(N5278), .Z(N5294) );
  CAN2X2 C41688 ( .A(N5266), .B(N5277), .Z(N5293) );
  CAN2X2 C41687 ( .A(N5266), .B(N5276), .Z(N5292) );
  CAN2X2 C41686 ( .A(N5266), .B(N5275), .Z(N5291) );
  CAN2X2 C41685 ( .A(N5266), .B(N5274), .Z(N5290) );
  CAN2X2 C41684 ( .A(N5266), .B(N5273), .Z(N5289) );
  CAN2X2 C41683 ( .A(N5265), .B(N5280), .Z(N5288) );
  CAN2X2 C41682 ( .A(N5265), .B(N5279), .Z(N5287) );
  CAN2X2 C41681 ( .A(N5265), .B(N5278), .Z(N5286) );
  CAN2X2 C41680 ( .A(N5265), .B(N5277), .Z(N5285) );
  CAN2X2 C41679 ( .A(N5265), .B(N5276), .Z(N5284) );
  CAN2X2 C41678 ( .A(N5265), .B(N5275), .Z(N5283) );
  CAN2X2 C41677 ( .A(N5265), .B(N5274), .Z(N5282) );
  CAN2X2 C41676 ( .A(N5265), .B(N5273), .Z(N5281) );
  CAN2X2 C41675 ( .A(N5124), .B(N5272), .Z(N5280) );
  CAN2X2 C41674 ( .A(N5124), .B(N5271), .Z(N5279) );
  CAN2X2 C41673 ( .A(N5124), .B(N5270), .Z(N5278) );
  CAN2X2 C41672 ( .A(N5124), .B(N5269), .Z(N5277) );
  CAN2X2 C41671 ( .A(write_ptr[2]), .B(N5272), .Z(N5276) );
  CAN2X2 C41670 ( .A(write_ptr[2]), .B(N5271), .Z(N5275) );
  CAN2X2 C41669 ( .A(write_ptr[2]), .B(N5270), .Z(N5274) );
  CAN2X2 C41668 ( .A(write_ptr[2]), .B(N5269), .Z(N5273) );
  CIVX2 I_35 ( .A(write_ptr[1]), .Z(N31) );
  CIVX2 I_34 ( .A(write_ptr[0]), .Z(N30) );
  CAN2X2 C41667 ( .A(N30), .B(N31), .Z(N5272) );
  CIVX2 I_33 ( .A(write_ptr[1]), .Z(N29) );
  CAN2X2 C41666 ( .A(write_ptr[0]), .B(N29), .Z(N5271) );
  CIVX2 I_32 ( .A(write_ptr[0]), .Z(N28) );
  CAN2X2 C41665 ( .A(N28), .B(write_ptr[1]), .Z(N5270) );
  CAN2X2 C41664 ( .A(write_ptr[0]), .B(write_ptr[1]), .Z(N5269) );
  CIVX2 I_31 ( .A(write_ptr[4]), .Z(N27) );
  CIVX2 I_30 ( .A(write_ptr[3]), .Z(N26) );
  CAN2X2 C41662 ( .A(N26), .B(N27), .Z(N5268) );
  CIVX2 I_29 ( .A(write_ptr[4]), .Z(N25) );
  CAN2X2 C41661 ( .A(write_ptr[3]), .B(N25), .Z(N5267) );
  CIVX2 I_28 ( .A(write_ptr[3]), .Z(N24) );
  CAN2X2 C41660 ( .A(N24), .B(write_ptr[4]), .Z(N5266) );
  CAN2X2 C41659 ( .A(write_ptr[3]), .B(write_ptr[4]), .Z(N5265) );
  CAN2X2 C41609 ( .A(N5220), .B(N5232), .Z(N5264) );
  CAN2X2 C41608 ( .A(N5220), .B(N5231), .Z(N5263) );
  CAN2X2 C41607 ( .A(N5220), .B(N5230), .Z(N5262) );
  CAN2X2 C41606 ( .A(N5220), .B(N5229), .Z(N5261) );
  CAN2X2 C41605 ( .A(N5220), .B(N5228), .Z(N5260) );
  CAN2X2 C41604 ( .A(N5220), .B(N5227), .Z(N5259) );
  CAN2X2 C41603 ( .A(N5220), .B(N5226), .Z(N5258) );
  CAN2X2 C41602 ( .A(N5220), .B(N5225), .Z(N5257) );
  CAN2X2 C41601 ( .A(N5219), .B(N5232), .Z(N5256) );
  CAN2X2 C41600 ( .A(N5219), .B(N5231), .Z(N5255) );
  CAN2X2 C41599 ( .A(N5219), .B(N5230), .Z(N5254) );
  CAN2X2 C41598 ( .A(N5219), .B(N5229), .Z(N5253) );
  CAN2X2 C41597 ( .A(N5219), .B(N5228), .Z(N5252) );
  CAN2X2 C41596 ( .A(N5219), .B(N5227), .Z(N5251) );
  CAN2X2 C41595 ( .A(N5219), .B(N5226), .Z(N5250) );
  CAN2X2 C41594 ( .A(N5219), .B(N5225), .Z(N5249) );
  CAN2X2 C41593 ( .A(N5218), .B(N5232), .Z(N5248) );
  CAN2X2 C41592 ( .A(N5218), .B(N5231), .Z(N5247) );
  CAN2X2 C41591 ( .A(N5218), .B(N5230), .Z(N5246) );
  CAN2X2 C41590 ( .A(N5218), .B(N5229), .Z(N5245) );
  CAN2X2 C41589 ( .A(N5218), .B(N5228), .Z(N5244) );
  CAN2X2 C41588 ( .A(N5218), .B(N5227), .Z(N5243) );
  CAN2X2 C41587 ( .A(N5218), .B(N5226), .Z(N5242) );
  CAN2X2 C41586 ( .A(N5218), .B(N5225), .Z(N5241) );
  CAN2X2 C41585 ( .A(N5217), .B(N5232), .Z(N5240) );
  CAN2X2 C41584 ( .A(N5217), .B(N5231), .Z(N5239) );
  CAN2X2 C41583 ( .A(N5217), .B(N5230), .Z(N5238) );
  CAN2X2 C41582 ( .A(N5217), .B(N5229), .Z(N5237) );
  CAN2X2 C41581 ( .A(N5217), .B(N5228), .Z(N5236) );
  CAN2X2 C41580 ( .A(N5217), .B(N5227), .Z(N5235) );
  CAN2X2 C41579 ( .A(N5217), .B(N5226), .Z(N5234) );
  CAN2X2 C41578 ( .A(N5217), .B(N5225), .Z(N5233) );
  CAN2X2 C41577 ( .A(N5124), .B(N5224), .Z(N5232) );
  CAN2X2 C41576 ( .A(N5124), .B(N5223), .Z(N5231) );
  CAN2X2 C41575 ( .A(N5124), .B(N5222), .Z(N5230) );
  CAN2X2 C41574 ( .A(N5124), .B(N5221), .Z(N5229) );
  CAN2X2 C41573 ( .A(write_ptr[2]), .B(N5224), .Z(N5228) );
  CAN2X2 C41572 ( .A(write_ptr[2]), .B(N5223), .Z(N5227) );
  CAN2X2 C41571 ( .A(write_ptr[2]), .B(N5222), .Z(N5226) );
  CAN2X2 C41570 ( .A(write_ptr[2]), .B(N5221), .Z(N5225) );
  CIVX2 I_27 ( .A(write_ptr[1]), .Z(N23) );
  CIVX2 I_26 ( .A(write_ptr[0]), .Z(N22) );
  CAN2X2 C41569 ( .A(N22), .B(N23), .Z(N5224) );
  CIVX2 I_25 ( .A(write_ptr[1]), .Z(N21) );
  CAN2X2 C41568 ( .A(write_ptr[0]), .B(N21), .Z(N5223) );
  CIVX2 I_24 ( .A(write_ptr[0]), .Z(N20) );
  CAN2X2 C41567 ( .A(N20), .B(write_ptr[1]), .Z(N5222) );
  CAN2X2 C41566 ( .A(write_ptr[0]), .B(write_ptr[1]), .Z(N5221) );
  CIVX2 I_23 ( .A(write_ptr[4]), .Z(N19) );
  CIVX2 I_22 ( .A(write_ptr[3]), .Z(N18) );
  CAN2X2 C41564 ( .A(N18), .B(N19), .Z(N5220) );
  CIVX2 I_21 ( .A(write_ptr[4]), .Z(N17) );
  CAN2X2 C41563 ( .A(write_ptr[3]), .B(N17), .Z(N5219) );
  CIVX2 I_20 ( .A(write_ptr[3]), .Z(N16) );
  CAN2X2 C41562 ( .A(N16), .B(write_ptr[4]), .Z(N5218) );
  CAN2X2 C41561 ( .A(write_ptr[3]), .B(write_ptr[4]), .Z(N5217) );
  CAN2X2 C41511 ( .A(N5172), .B(N5184), .Z(N5216) );
  CAN2X2 C41510 ( .A(N5172), .B(N5183), .Z(N5215) );
  CAN2X2 C41509 ( .A(N5172), .B(N5182), .Z(N5214) );
  CAN2X2 C41508 ( .A(N5172), .B(N5181), .Z(N5213) );
  CAN2X2 C41507 ( .A(N5172), .B(N5180), .Z(N5212) );
  CAN2X2 C41506 ( .A(N5172), .B(N5179), .Z(N5211) );
  CAN2X2 C41505 ( .A(N5172), .B(N5178), .Z(N5210) );
  CAN2X2 C41504 ( .A(N5172), .B(N5177), .Z(N5209) );
  CAN2X2 C41503 ( .A(N5171), .B(N5184), .Z(N5208) );
  CAN2X2 C41502 ( .A(N5171), .B(N5183), .Z(N5207) );
  CAN2X2 C41501 ( .A(N5171), .B(N5182), .Z(N5206) );
  CAN2X2 C41500 ( .A(N5171), .B(N5181), .Z(N5205) );
  CAN2X2 C41499 ( .A(N5171), .B(N5180), .Z(N5204) );
  CAN2X2 C41498 ( .A(N5171), .B(N5179), .Z(N5203) );
  CAN2X2 C41497 ( .A(N5171), .B(N5178), .Z(N5202) );
  CAN2X2 C41496 ( .A(N5171), .B(N5177), .Z(N5201) );
  CAN2X2 C41495 ( .A(N5170), .B(N5184), .Z(N5200) );
  CAN2X2 C41494 ( .A(N5170), .B(N5183), .Z(N5199) );
  CAN2X2 C41493 ( .A(N5170), .B(N5182), .Z(N5198) );
  CAN2X2 C41492 ( .A(N5170), .B(N5181), .Z(N5197) );
  CAN2X2 C41491 ( .A(N5170), .B(N5180), .Z(N5196) );
  CAN2X2 C41490 ( .A(N5170), .B(N5179), .Z(N5195) );
  CAN2X2 C41489 ( .A(N5170), .B(N5178), .Z(N5194) );
  CAN2X2 C41488 ( .A(N5170), .B(N5177), .Z(N5193) );
  CAN2X2 C41487 ( .A(N5169), .B(N5184), .Z(N5192) );
  CAN2X2 C41486 ( .A(N5169), .B(N5183), .Z(N5191) );
  CAN2X2 C41485 ( .A(N5169), .B(N5182), .Z(N5190) );
  CAN2X2 C41484 ( .A(N5169), .B(N5181), .Z(N5189) );
  CAN2X2 C41483 ( .A(N5169), .B(N5180), .Z(N5188) );
  CAN2X2 C41482 ( .A(N5169), .B(N5179), .Z(N5187) );
  CAN2X2 C41481 ( .A(N5169), .B(N5178), .Z(N5186) );
  CAN2X2 C41480 ( .A(N5169), .B(N5177), .Z(N5185) );
  CAN2X2 C41479 ( .A(N5124), .B(N5176), .Z(N5184) );
  CAN2X2 C41478 ( .A(N5124), .B(N5175), .Z(N5183) );
  CAN2X2 C41477 ( .A(N5124), .B(N5174), .Z(N5182) );
  CAN2X2 C41476 ( .A(N5124), .B(N5173), .Z(N5181) );
  CAN2X2 C41475 ( .A(write_ptr[2]), .B(N5176), .Z(N5180) );
  CAN2X2 C41474 ( .A(write_ptr[2]), .B(N5175), .Z(N5179) );
  CAN2X2 C41473 ( .A(write_ptr[2]), .B(N5174), .Z(N5178) );
  CAN2X2 C41472 ( .A(write_ptr[2]), .B(N5173), .Z(N5177) );
  CIVX2 I_19 ( .A(write_ptr[1]), .Z(N15) );
  CIVX2 I_18 ( .A(write_ptr[0]), .Z(N14) );
  CAN2X2 C41471 ( .A(N14), .B(N15), .Z(N5176) );
  CIVX2 I_17 ( .A(write_ptr[1]), .Z(N13) );
  CAN2X2 C41470 ( .A(write_ptr[0]), .B(N13), .Z(N5175) );
  CIVX2 I_16 ( .A(write_ptr[0]), .Z(N12) );
  CAN2X2 C41469 ( .A(N12), .B(write_ptr[1]), .Z(N5174) );
  CAN2X2 C41468 ( .A(write_ptr[0]), .B(write_ptr[1]), .Z(N5173) );
  CIVX2 I_15 ( .A(write_ptr[4]), .Z(N11) );
  CIVX2 I_14 ( .A(write_ptr[3]), .Z(N10) );
  CAN2X2 C41466 ( .A(N10), .B(N11), .Z(N5172) );
  CIVX2 I_13 ( .A(write_ptr[4]), .Z(N9) );
  CAN2X2 C41465 ( .A(write_ptr[3]), .B(N9), .Z(N5171) );
  CIVX2 I_12 ( .A(write_ptr[3]), .Z(N8) );
  CAN2X2 C41464 ( .A(N8), .B(write_ptr[4]), .Z(N5170) );
  CAN2X2 C41463 ( .A(write_ptr[3]), .B(write_ptr[4]), .Z(N5169) );
  CAN2X2 C41413 ( .A(N5123), .B(N5136), .Z(N5168) );
  CAN2X2 C41412 ( .A(N5123), .B(N5135), .Z(N5167) );
  CAN2X2 C41411 ( .A(N5123), .B(N5134), .Z(N5166) );
  CAN2X2 C41410 ( .A(N5123), .B(N5133), .Z(N5165) );
  CAN2X2 C41409 ( .A(N5123), .B(N5132), .Z(N5164) );
  CAN2X2 C41408 ( .A(N5123), .B(N5131), .Z(N5163) );
  CAN2X2 C41407 ( .A(N5123), .B(N5130), .Z(N5162) );
  CAN2X2 C41406 ( .A(N5123), .B(N5129), .Z(N5161) );
  CAN2X2 C41405 ( .A(N5122), .B(N5136), .Z(N5160) );
  CAN2X2 C41404 ( .A(N5122), .B(N5135), .Z(N5159) );
  CAN2X2 C41403 ( .A(N5122), .B(N5134), .Z(N5158) );
  CAN2X2 C41402 ( .A(N5122), .B(N5133), .Z(N5157) );
  CAN2X2 C41401 ( .A(N5122), .B(N5132), .Z(N5156) );
  CAN2X2 C41400 ( .A(N5122), .B(N5131), .Z(N5155) );
  CAN2X2 C41399 ( .A(N5122), .B(N5130), .Z(N5154) );
  CAN2X2 C41398 ( .A(N5122), .B(N5129), .Z(N5153) );
  CAN2X2 C41397 ( .A(N5121), .B(N5136), .Z(N5152) );
  CAN2X2 C41396 ( .A(N5121), .B(N5135), .Z(N5151) );
  CAN2X2 C41395 ( .A(N5121), .B(N5134), .Z(N5150) );
  CAN2X2 C41394 ( .A(N5121), .B(N5133), .Z(N5149) );
  CAN2X2 C41393 ( .A(N5121), .B(N5132), .Z(N5148) );
  CAN2X2 C41392 ( .A(N5121), .B(N5131), .Z(N5147) );
  CAN2X2 C41391 ( .A(N5121), .B(N5130), .Z(N5146) );
  CAN2X2 C41390 ( .A(N5121), .B(N5129), .Z(N5145) );
  CAN2X2 C41389 ( .A(N5120), .B(N5136), .Z(N5144) );
  CAN2X2 C41388 ( .A(N5120), .B(N5135), .Z(N5143) );
  CAN2X2 C41387 ( .A(N5120), .B(N5134), .Z(N5142) );
  CAN2X2 C41386 ( .A(N5120), .B(N5133), .Z(N5141) );
  CAN2X2 C41385 ( .A(N5120), .B(N5132), .Z(N5140) );
  CAN2X2 C41384 ( .A(N5120), .B(N5131), .Z(N5139) );
  CAN2X2 C41383 ( .A(N5120), .B(N5130), .Z(N5138) );
  CAN2X2 C41382 ( .A(N5120), .B(N5129), .Z(N5137) );
  CAN2X2 C41381 ( .A(N5124), .B(N5128), .Z(N5136) );
  CAN2X2 C41380 ( .A(N5124), .B(N5127), .Z(N5135) );
  CAN2X2 C41379 ( .A(N5124), .B(N5126), .Z(N5134) );
  CAN2X2 C41378 ( .A(N5124), .B(N5125), .Z(N5133) );
  CAN2X2 C41377 ( .A(write_ptr[2]), .B(N5128), .Z(N5132) );
  CAN2X2 C41376 ( .A(write_ptr[2]), .B(N5127), .Z(N5131) );
  CAN2X2 C41375 ( .A(write_ptr[2]), .B(N5126), .Z(N5130) );
  CAN2X2 C41374 ( .A(write_ptr[2]), .B(N5125), .Z(N5129) );
  CIVX2 I_11 ( .A(write_ptr[1]), .Z(N7) );
  CIVX2 I_10 ( .A(write_ptr[0]), .Z(N6) );
  CAN2X2 C41373 ( .A(N6), .B(N7), .Z(N5128) );
  CIVX2 I_9 ( .A(write_ptr[1]), .Z(N5) );
  CAN2X2 C41372 ( .A(write_ptr[0]), .B(N5), .Z(N5127) );
  CIVX2 I_8 ( .A(write_ptr[0]), .Z(N4) );
  CAN2X2 C41371 ( .A(N4), .B(write_ptr[1]), .Z(N5126) );
  CAN2X2 C41370 ( .A(write_ptr[0]), .B(write_ptr[1]), .Z(N5125) );
  CIVX2 I_7 ( .A(write_ptr[2]), .Z(N5124) );
  CIVX2 I_6 ( .A(write_ptr[4]), .Z(N3) );
  CIVX2 I_5 ( .A(write_ptr[3]), .Z(N2) );
  CAN2X2 C41368 ( .A(N2), .B(N3), .Z(N5123) );
  CIVX2 I_4 ( .A(write_ptr[4]), .Z(N1) );
  CAN2X2 C41367 ( .A(write_ptr[3]), .B(N1), .Z(N5122) );
  CIVX2 I_3 ( .A(write_ptr[3]), .Z(N0) );
  CAN2X2 C41366 ( .A(N0), .B(write_ptr[4]), .Z(N5121) );
  CAN2X2 C41365 ( .A(write_ptr[3]), .B(write_ptr[4]), .Z(N5120) );
  COR3X1 C36753 ( .A(N210), .B(N4965), .C(N213), .Z(N2531) );
  COR3X1 C36530 ( .A(N210), .B(n2610), .C(N213), .Z(N2525) );
  CIVX2 I_2 ( .A(N5117), .Z(N5118) );
  COR2X1 C36454 ( .A(counter[0]), .B(N5116), .Z(N5117) );
  COR2X1 C36453 ( .A(counter[1]), .B(N5115), .Z(N5116) );
  COR2X1 C36452 ( .A(counter[2]), .B(N5114), .Z(N5115) );
  COR2X1 C36451 ( .A(counter[3]), .B(N5113), .Z(N5114) );
  CIVX2 I_1 ( .A(N5111), .Z(N5112) );
  COR2X1 C36448 ( .A(counter[0]), .B(N5110), .Z(N5111) );
  COR2X1 C36447 ( .A(counter[1]), .B(N5109), .Z(N5110) );
  COR2X1 C36446 ( .A(counter[2]), .B(N5108), .Z(N5109) );
  COR2X1 C36445 ( .A(counter[3]), .B(N5107), .Z(N5108) );
  CFD2QX1 \out_reg[0]  ( .D(n2529), .CP(clk), .CD(n77), .Q(out[0]) );
  CFD2QX1 \out_reg[1]  ( .D(n2528), .CP(clk), .CD(n77), .Q(out[1]) );
  CFD2QX1 \out_reg[2]  ( .D(n2527), .CP(clk), .CD(n77), .Q(out[2]) );
  CFD2QX1 \out_reg[3]  ( .D(n2526), .CP(clk), .CD(n77), .Q(out[3]) );
  CFD2QX1 \out_reg[4]  ( .D(n2525), .CP(clk), .CD(n77), .Q(out[4]) );
  CFD2QX1 \out_reg[5]  ( .D(n2524), .CP(clk), .CD(n77), .Q(out[5]) );
  CFD2QX1 \out_reg[6]  ( .D(n2523), .CP(clk), .CD(n77), .Q(out[6]) );
  CFD2QX1 \out_reg[7]  ( .D(n2522), .CP(clk), .CD(n77), .Q(out[7]) );
  CFD2QX1 \out_reg[8]  ( .D(n2521), .CP(clk), .CD(n77), .Q(out[8]) );
  CFD2QX1 \out_reg[9]  ( .D(n2520), .CP(clk), .CD(n77), .Q(out[9]) );
  CFD2QX1 \out_reg[10]  ( .D(n2519), .CP(clk), .CD(n77), .Q(out[10]) );
  CFD2QX1 \out_reg[11]  ( .D(n2518), .CP(clk), .CD(n77), .Q(out[11]) );
  CFD2QX1 \out_reg[12]  ( .D(n2517), .CP(clk), .CD(n77), .Q(out[12]) );
  CFD2QX1 \out_reg[13]  ( .D(n2516), .CP(clk), .CD(n77), .Q(out[13]) );
  CFD2QX1 \out_reg[14]  ( .D(n2515), .CP(clk), .CD(n77), .Q(out[14]) );
  CFD2QX1 \out_reg[15]  ( .D(n2514), .CP(clk), .CD(n77), .Q(out[15]) );
  CFD2QX1 \out_reg[16]  ( .D(n2513), .CP(clk), .CD(n77), .Q(out[16]) );
  CFD2QX1 \out_reg[17]  ( .D(n2512), .CP(clk), .CD(n77), .Q(out[17]) );
  CFD2QX1 \out_reg[18]  ( .D(n2511), .CP(clk), .CD(n77), .Q(out[18]) );
  CFD2QX1 \out_reg[19]  ( .D(n2510), .CP(clk), .CD(n77), .Q(out[19]) );
  CFD2QX1 \out_reg[20]  ( .D(n2509), .CP(clk), .CD(n77), .Q(out[20]) );
  CFD2QX1 \out_reg[21]  ( .D(n2508), .CP(clk), .CD(n77), .Q(out[21]) );
  CFD2QX1 \out_reg[22]  ( .D(n2507), .CP(clk), .CD(n77), .Q(out[22]) );
  CFD2QX1 \out_reg[23]  ( .D(n2506), .CP(clk), .CD(n77), .Q(out[23]) );
  CFD2QX1 \out_reg[24]  ( .D(n2505), .CP(clk), .CD(n77), .Q(out[24]) );
  CFD2QX1 \out_reg[25]  ( .D(n2504), .CP(clk), .CD(n77), .Q(out[25]) );
  CFD2QX1 \out_reg[26]  ( .D(n2503), .CP(clk), .CD(n77), .Q(out[26]) );
  CFD2QX1 \out_reg[27]  ( .D(n2502), .CP(clk), .CD(n77), .Q(out[27]) );
  CFD2QX1 \out_reg[28]  ( .D(n2501), .CP(clk), .CD(n77), .Q(out[28]) );
  CFD2QX1 \out_reg[29]  ( .D(n2500), .CP(clk), .CD(n77), .Q(out[29]) );
  CFD2QX1 \out_reg[30]  ( .D(n2499), .CP(clk), .CD(n77), .Q(out[30]) );
  CFD2QX1 \out_reg[31]  ( .D(n2498), .CP(clk), .CD(n77), .Q(out[31]) );
  CFD2QX1 \out_reg[32]  ( .D(n2497), .CP(clk), .CD(n77), .Q(out[32]) );
  CFD2QX1 \out_reg[33]  ( .D(n2496), .CP(clk), .CD(n77), .Q(out[33]) );
  CFD2QX1 \out_reg[34]  ( .D(n2495), .CP(clk), .CD(n77), .Q(out[34]) );
  CFD2QX1 \out_reg[35]  ( .D(n2494), .CP(clk), .CD(n77), .Q(out[35]) );
  CFD2QX1 \out_reg[36]  ( .D(n2493), .CP(clk), .CD(n77), .Q(out[36]) );
  CFD2QX1 \out_reg[37]  ( .D(n2492), .CP(clk), .CD(n77), .Q(out[37]) );
  CFD2QX1 \out_reg[38]  ( .D(n2491), .CP(clk), .CD(n77), .Q(out[38]) );
  CFD2QX1 \out_reg[39]  ( .D(n2490), .CP(clk), .CD(n77), .Q(out[39]) );
  CFD2QX1 \out_reg[40]  ( .D(n2489), .CP(clk), .CD(n77), .Q(out[40]) );
  CFD2QX1 \out_reg[41]  ( .D(n2488), .CP(clk), .CD(n77), .Q(out[41]) );
  CFD2QX1 \out_reg[42]  ( .D(n2487), .CP(clk), .CD(n77), .Q(out[42]) );
  CFD2QX1 \out_reg[43]  ( .D(n2486), .CP(clk), .CD(n77), .Q(out[43]) );
  CFD2QX1 \out_reg[44]  ( .D(n2485), .CP(clk), .CD(n77), .Q(out[44]) );
  CFD2QX1 \out_reg[45]  ( .D(n2484), .CP(clk), .CD(n77), .Q(out[45]) );
  CFD2QX1 \out_reg[46]  ( .D(n2483), .CP(clk), .CD(n77), .Q(out[46]) );
  CFD2QX1 \out_reg[47]  ( .D(n2482), .CP(clk), .CD(n77), .Q(out[47]) );
  CFD2QX1 \out_reg[48]  ( .D(n2481), .CP(clk), .CD(n77), .Q(out[48]) );
  CFD2QX1 \out_reg[49]  ( .D(n2480), .CP(clk), .CD(n77), .Q(out[49]) );
  CFD2QX1 \out_reg[50]  ( .D(n2479), .CP(clk), .CD(n77), .Q(out[50]) );
  CFD2QX1 \out_reg[51]  ( .D(n2478), .CP(clk), .CD(n77), .Q(out[51]) );
  CFD2QX1 \out_reg[52]  ( .D(n2477), .CP(clk), .CD(n77), .Q(out[52]) );
  CFD2QX1 \out_reg[53]  ( .D(n2476), .CP(clk), .CD(n77), .Q(out[53]) );
  CFD2QX1 \out_reg[54]  ( .D(n2475), .CP(clk), .CD(n77), .Q(out[54]) );
  CFD2QX1 \out_reg[55]  ( .D(n2474), .CP(clk), .CD(n77), .Q(out[55]) );
  CFD2QX1 \out_reg[56]  ( .D(n2473), .CP(clk), .CD(n77), .Q(out[56]) );
  CFD2QX1 \out_reg[57]  ( .D(n2472), .CP(clk), .CD(n77), .Q(out[57]) );
  CFD2QX1 \out_reg[58]  ( .D(n2471), .CP(clk), .CD(n77), .Q(out[58]) );
  CFD2QX1 \out_reg[59]  ( .D(n2470), .CP(clk), .CD(n77), .Q(out[59]) );
  CFD2QX1 \out_reg[60]  ( .D(n2469), .CP(clk), .CD(n77), .Q(out[60]) );
  CFD2QX1 \out_reg[61]  ( .D(n2468), .CP(clk), .CD(n77), .Q(out[61]) );
  CFD2QX1 \out_reg[62]  ( .D(n2467), .CP(clk), .CD(n77), .Q(out[62]) );
  CFD2QX1 \lout_reg[0]  ( .D(n2466), .CP(clk), .CD(n77), .Q(lout[0]) );
  CFD2QX1 \lout_reg[1]  ( .D(n2535), .CP(clk), .CD(n77), .Q(lout[1]) );
  CFD2QX1 \lout_reg[2]  ( .D(n2534), .CP(clk), .CD(n77), .Q(lout[2]) );
  CFD2QX1 \lout_reg[3]  ( .D(n2533), .CP(clk), .CD(n77), .Q(lout[3]) );
  CFD2QX1 \lout_reg[4]  ( .D(n2532), .CP(clk), .CD(n77), .Q(lout[4]) );
  CFD2QX1 \lout_reg[5]  ( .D(n2531), .CP(clk), .CD(n77), .Q(lout[5]) );
  CFD2QX1 \lout_reg[6]  ( .D(n2530), .CP(clk), .CD(n77), .Q(lout[6]) );
  CFD2QX1 \counter_reg[0]  ( .D(n2459), .CP(clk), .CD(n77), .Q(counter[0]) );
  CFD2X1 \counter_reg[5]  ( .D(n2458), .CP(clk), .CD(n77), .Q(counter[5]), 
        .QN(N5106) );
  CFD2QX1 \counter_reg[1]  ( .D(n2454), .CP(clk), .CD(n77), .Q(counter[1]) );
  CFD2QX1 \counter_reg[4]  ( .D(n2457), .CP(clk), .CD(n77), .Q(counter[4]) );
  CFD2QX1 \counter_reg[2]  ( .D(n2455), .CP(clk), .CD(n77), .Q(counter[2]) );
  CFD2QX1 \counter_reg[3]  ( .D(n2456), .CP(clk), .CD(n77), .Q(counter[3]) );
  CFD2QX1 \read_ptr_reg[0]  ( .D(n2382), .CP(clk), .CD(n77), .Q(N38) );
  CFD2QX1 \read_ptr_reg[1]  ( .D(n2381), .CP(clk), .CD(n77), .Q(N39) );
  CFD2QX1 \read_ptr_reg[2]  ( .D(n2380), .CP(clk), .CD(n77), .Q(N40) );
  CFD2QX1 \write_ptr_reg[0]  ( .D(n2377), .CP(clk), .CD(n77), .Q(write_ptr[0])
         );
  CFD2QX1 \write_ptr_reg[1]  ( .D(n2376), .CP(clk), .CD(n77), .Q(write_ptr[1])
         );
  CFD2QX1 \write_ptr_reg[2]  ( .D(n2375), .CP(clk), .CD(n77), .Q(write_ptr[2])
         );
  CFD2QX1 \write_ptr_reg[3]  ( .D(n2374), .CP(clk), .CD(n77), .Q(write_ptr[3])
         );
  CFD2QX1 \write_ptr_reg[4]  ( .D(n2373), .CP(clk), .CD(n77), .Q(write_ptr[4])
         );
  CAOR2X1 U3 ( .A(N132), .B(n2), .C(lout_new[6]), .D(n3), .Z(n6) );
  CAOR2X1 U4 ( .A(N131), .B(n2), .C(lout_new[5]), .D(n3), .Z(n7) );
  CAOR2X1 U5 ( .A(N130), .B(n2), .C(lout_new[4]), .D(n3), .Z(n8) );
  CAOR2X1 U6 ( .A(N129), .B(n2), .C(lout_new[3]), .D(n3), .Z(n9) );
  CAOR2X1 U7 ( .A(N128), .B(n2), .C(lout_new[2]), .D(n3), .Z(n10) );
  CAOR2X1 U8 ( .A(N127), .B(n2), .C(lout_new[1]), .D(n3), .Z(n11) );
  CAOR2X1 U9 ( .A(N126), .B(n2), .C(lout_new[0]), .D(n3), .Z(n12) );
  CAOR2X1 U10 ( .A(datain), .B(n2), .C(out_new[0]), .D(n3), .Z(n13) );
  CAOR2X1 U11 ( .A(n2598), .B(n2), .C(out_new[1]), .D(n3), .Z(n14) );
  CAOR2X1 U12 ( .A(n2597), .B(n2), .C(out_new[2]), .D(n3), .Z(n15) );
  CAOR2X1 U13 ( .A(n2596), .B(n2), .C(out_new[3]), .D(n3), .Z(n16) );
  CAOR2X1 U14 ( .A(n2595), .B(n2), .C(out_new[4]), .D(n3), .Z(n17) );
  CAOR2X1 U15 ( .A(n2594), .B(n2), .C(out_new[5]), .D(n3), .Z(n18) );
  CAOR2X1 U16 ( .A(n2593), .B(n2), .C(out_new[6]), .D(n3), .Z(n19) );
  CAOR2X1 U17 ( .A(n2592), .B(n2), .C(out_new[7]), .D(n3), .Z(n20) );
  CAOR2X1 U18 ( .A(n2591), .B(n2), .C(out_new[8]), .D(n3), .Z(n21) );
  CAOR2X1 U19 ( .A(n2590), .B(n2), .C(out_new[9]), .D(n3), .Z(n22) );
  CAOR2X1 U20 ( .A(n2589), .B(n2), .C(out_new[10]), .D(n3), .Z(n23) );
  CAOR2X1 U21 ( .A(n2588), .B(n2), .C(out_new[11]), .D(n3), .Z(n24) );
  CAOR2X1 U22 ( .A(n2587), .B(n2), .C(out_new[12]), .D(n3), .Z(n25) );
  CAOR2X1 U23 ( .A(n2586), .B(n2), .C(out_new[13]), .D(n3), .Z(n26) );
  CAOR2X1 U24 ( .A(n2585), .B(n2), .C(out_new[14]), .D(n3), .Z(n27) );
  CAOR2X1 U25 ( .A(n2584), .B(n2), .C(out_new[15]), .D(n3), .Z(n28) );
  CAOR2X1 U26 ( .A(n2583), .B(n2), .C(out_new[16]), .D(n3), .Z(n29) );
  CAOR2X1 U27 ( .A(n2582), .B(n2), .C(out_new[17]), .D(n3), .Z(n30) );
  CAOR2X1 U28 ( .A(n2581), .B(n2), .C(out_new[18]), .D(n3), .Z(n31) );
  CAOR2X1 U29 ( .A(n2580), .B(n2), .C(out_new[19]), .D(n3), .Z(n32) );
  CAOR2X1 U30 ( .A(n2579), .B(n2), .C(out_new[20]), .D(n3), .Z(n33) );
  CAOR2X1 U31 ( .A(n2578), .B(n2), .C(out_new[21]), .D(n3), .Z(n34) );
  CAOR2X1 U32 ( .A(n2577), .B(n2), .C(out_new[22]), .D(n3), .Z(n35) );
  CAOR2X1 U33 ( .A(n2576), .B(n2), .C(out_new[23]), .D(n3), .Z(n36) );
  CAOR2X1 U34 ( .A(n2575), .B(n2), .C(out_new[24]), .D(n3), .Z(n37) );
  CAOR2X1 U35 ( .A(n2574), .B(n2), .C(out_new[25]), .D(n3), .Z(n38) );
  CAOR2X1 U36 ( .A(n2573), .B(n2), .C(out_new[26]), .D(n3), .Z(n39) );
  CAOR2X1 U37 ( .A(n2572), .B(n2), .C(out_new[27]), .D(n3), .Z(n40) );
  CAOR2X1 U38 ( .A(n2571), .B(n2), .C(out_new[28]), .D(n3), .Z(n41) );
  CAOR2X1 U39 ( .A(n2570), .B(n2), .C(out_new[29]), .D(n3), .Z(n42) );
  CAOR2X1 U40 ( .A(n2569), .B(n2), .C(out_new[30]), .D(n3), .Z(n43) );
  CAOR2X1 U41 ( .A(n2568), .B(n2), .C(out_new[31]), .D(n3), .Z(n44) );
  CAOR2X1 U42 ( .A(n2567), .B(n2), .C(out_new[32]), .D(n3), .Z(n45) );
  CAOR2X1 U43 ( .A(n2566), .B(n2), .C(out_new[33]), .D(n3), .Z(n46) );
  CAOR2X1 U44 ( .A(n2565), .B(n2), .C(out_new[34]), .D(n3), .Z(n47) );
  CAOR2X1 U45 ( .A(n2564), .B(n2), .C(out_new[35]), .D(n3), .Z(n48) );
  CAOR2X1 U46 ( .A(n2563), .B(n2), .C(out_new[36]), .D(n3), .Z(n49) );
  CAOR2X1 U47 ( .A(n2562), .B(n2), .C(out_new[37]), .D(n3), .Z(n50) );
  CAOR2X1 U48 ( .A(n2561), .B(n2), .C(out_new[38]), .D(n3), .Z(n51) );
  CAOR2X1 U49 ( .A(n2560), .B(n2), .C(out_new[39]), .D(n3), .Z(n52) );
  CAOR2X1 U50 ( .A(n2559), .B(n2), .C(out_new[40]), .D(n3), .Z(n53) );
  CAOR2X1 U51 ( .A(n2558), .B(n2), .C(out_new[41]), .D(n3), .Z(n54) );
  CAOR2X1 U52 ( .A(n2557), .B(n2), .C(out_new[42]), .D(n3), .Z(n55) );
  CAOR2X1 U53 ( .A(n2556), .B(n2), .C(out_new[43]), .D(n3), .Z(n56) );
  CAOR2X1 U54 ( .A(n2555), .B(n2), .C(out_new[44]), .D(n3), .Z(n57) );
  CAOR2X1 U55 ( .A(n2554), .B(n2), .C(out_new[45]), .D(n3), .Z(n58) );
  CAOR2X1 U56 ( .A(n2553), .B(n2), .C(out_new[46]), .D(n3), .Z(n59) );
  CAOR2X1 U57 ( .A(n2552), .B(n2), .C(out_new[47]), .D(n3), .Z(n60) );
  CAOR2X1 U58 ( .A(n2551), .B(n2), .C(out_new[48]), .D(n3), .Z(n61) );
  CAOR2X1 U59 ( .A(n2550), .B(n2), .C(out_new[49]), .D(n3), .Z(n62) );
  CAOR2X1 U60 ( .A(n2549), .B(n2), .C(out_new[50]), .D(n3), .Z(n63) );
  CAOR2X1 U61 ( .A(n2548), .B(n2), .C(out_new[51]), .D(n3), .Z(n64) );
  CAOR2X1 U62 ( .A(n2547), .B(n2), .C(out_new[52]), .D(n3), .Z(n65) );
  CAOR2X1 U63 ( .A(n2546), .B(n2), .C(out_new[53]), .D(n3), .Z(n66) );
  CAOR2X1 U64 ( .A(n2545), .B(n2), .C(out_new[54]), .D(n3), .Z(n67) );
  CAOR2X1 U65 ( .A(n2544), .B(n2), .C(out_new[55]), .D(n3), .Z(n68) );
  CAOR2X1 U66 ( .A(n2543), .B(n2), .C(out_new[56]), .D(n3), .Z(n69) );
  CAOR2X1 U67 ( .A(n2542), .B(n2), .C(out_new[57]), .D(n3), .Z(n70) );
  CAOR2X1 U68 ( .A(n2541), .B(n2), .C(out_new[58]), .D(n3), .Z(n71) );
  CAOR2X1 U69 ( .A(n2540), .B(n2), .C(out_new[59]), .D(n3), .Z(n72) );
  CAOR2X1 U70 ( .A(n2539), .B(n2), .C(out_new[60]), .D(n3), .Z(n73) );
  CAOR2X1 U71 ( .A(n2538), .B(n2), .C(out_new[61]), .D(n3), .Z(n74) );
  CAOR2X1 U72 ( .A(n2537), .B(n2), .C(out_new[62]), .D(n3), .Z(n75) );
  CAOR2X1 U73 ( .A(n2536), .B(n2), .C(out_new[63]), .D(n3), .Z(n76) );
  CIVX1 U74 ( .A(n3), .Z(n2) );
  CNR2X1 U76 ( .A(n78), .B(n79), .Z(N123) );
  CIVX1 U82 ( .A(n80), .Z(N4965) );
  CAOR2X1 U85 ( .A(N5185), .B(n82), .C(N5281), .D(n83), .Z(N4818) );
  CAOR2X1 U87 ( .A(N5186), .B(n82), .C(N5282), .D(n83), .Z(N4747) );
  CAOR2X1 U89 ( .A(N5187), .B(n82), .C(N5283), .D(n83), .Z(N4676) );
  CAOR2X1 U91 ( .A(N5188), .B(n82), .C(N5284), .D(n83), .Z(N4605) );
  CAOR2X1 U93 ( .A(N5189), .B(n82), .C(N5285), .D(n83), .Z(N4534) );
  CAOR2X1 U95 ( .A(N5190), .B(n82), .C(N5286), .D(n83), .Z(N4463) );
  CAOR2X1 U97 ( .A(N5191), .B(n82), .C(N5287), .D(n83), .Z(N4392) );
  CAOR2X1 U99 ( .A(N5192), .B(n82), .C(N5288), .D(n83), .Z(N4321) );
  CAOR2X1 U101 ( .A(N5193), .B(n82), .C(N5289), .D(n83), .Z(N4250) );
  CAOR2X1 U103 ( .A(N5194), .B(n82), .C(N5290), .D(n83), .Z(N4179) );
  CAOR2X1 U105 ( .A(N5195), .B(n82), .C(N5291), .D(n83), .Z(N4108) );
  CAOR2X1 U107 ( .A(N5196), .B(n82), .C(N5292), .D(n83), .Z(N4037) );
  CAOR2X1 U109 ( .A(N5197), .B(n82), .C(N5293), .D(n83), .Z(N3966) );
  CAOR2X1 U111 ( .A(N5198), .B(n82), .C(N5294), .D(n83), .Z(N3895) );
  CAOR2X1 U113 ( .A(N5199), .B(n82), .C(N5295), .D(n83), .Z(N3824) );
  CAOR2X1 U115 ( .A(N5200), .B(n82), .C(N5296), .D(n83), .Z(N3753) );
  CAOR2X1 U117 ( .A(N5201), .B(n82), .C(N5297), .D(n83), .Z(N3682) );
  CAOR2X1 U119 ( .A(N5202), .B(n82), .C(N5298), .D(n83), .Z(N3611) );
  CAOR2X1 U121 ( .A(N5203), .B(n82), .C(N5299), .D(n83), .Z(N3540) );
  CAOR2X1 U123 ( .A(N5204), .B(n82), .C(N5300), .D(n83), .Z(N3469) );
  CAOR2X1 U125 ( .A(N5205), .B(n82), .C(N5301), .D(n83), .Z(N3398) );
  CAOR2X1 U127 ( .A(N5206), .B(n82), .C(N5302), .D(n83), .Z(N3327) );
  CAOR2X1 U129 ( .A(N5207), .B(n82), .C(N5303), .D(n83), .Z(N3256) );
  CAOR2X1 U131 ( .A(N5208), .B(n82), .C(N5304), .D(n83), .Z(N3185) );
  CAOR2X1 U133 ( .A(N5209), .B(n82), .C(N5305), .D(n83), .Z(N3114) );
  CAOR2X1 U135 ( .A(N5210), .B(n82), .C(N5306), .D(n83), .Z(N3043) );
  CAOR2X1 U137 ( .A(N5211), .B(n82), .C(N5307), .D(n83), .Z(N2972) );
  CAOR2X1 U139 ( .A(N5212), .B(n82), .C(N5308), .D(n83), .Z(N2901) );
  CAOR2X1 U141 ( .A(N5213), .B(n82), .C(N5309), .D(n83), .Z(N2830) );
  CAOR2X1 U143 ( .A(N5214), .B(n82), .C(N5310), .D(n83), .Z(N2759) );
  CAOR2X1 U145 ( .A(N5215), .B(n82), .C(N5311), .D(n83), .Z(N2688) );
  CAOR2X1 U147 ( .A(N5216), .B(n82), .C(N5312), .D(n83), .Z(N2617) );
  CND2X1 U152 ( .A(N235), .B(N114), .Z(n86) );
  CND2X1 U153 ( .A(N247), .B(n87), .Z(n85) );
  CND2X1 U154 ( .A(n88), .B(n89), .Z(N2537) );
  CND2X1 U155 ( .A(N234), .B(N114), .Z(n89) );
  CND2X1 U157 ( .A(n91), .B(n92), .Z(N2536) );
  CND2X1 U158 ( .A(N233), .B(N114), .Z(n92) );
  CANR2X1 U159 ( .A(counter[3]), .B(n90), .C(N245), .D(n87), .Z(n91) );
  CND2X1 U160 ( .A(n93), .B(n94), .Z(N2535) );
  CND2X1 U161 ( .A(N232), .B(N114), .Z(n94) );
  CANR2X1 U162 ( .A(counter[2]), .B(n90), .C(N244), .D(n87), .Z(n93) );
  CND2X1 U163 ( .A(n95), .B(n96), .Z(N2534) );
  CND2X1 U164 ( .A(N231), .B(N114), .Z(n96) );
  CANR2X1 U165 ( .A(counter[1]), .B(n90), .C(N243), .D(n87), .Z(n95) );
  CND2X1 U166 ( .A(n97), .B(n98), .Z(N2533) );
  CND2X1 U167 ( .A(N230), .B(N114), .Z(n98) );
  CANR2X1 U168 ( .A(counter[0]), .B(n90), .C(N242), .D(n87), .Z(n97) );
  CAOR2X1 U169 ( .A(N42), .B(N213), .C(N223), .D(n99), .Z(N2532) );
  CAOR2X1 U170 ( .A(N41), .B(N213), .C(N222), .D(n99), .Z(N2530) );
  CAOR2X1 U171 ( .A(n2623), .B(N213), .C(N221), .D(n99), .Z(N2529) );
  CAOR2X1 U172 ( .A(n2635), .B(N213), .C(N220), .D(n99), .Z(N2528) );
  CAOR2X1 U173 ( .A(n2647), .B(N213), .C(n2648), .D(n99), .Z(N2527) );
  CND2X1 U174 ( .A(N4961), .B(n80), .Z(n99) );
  CND2X1 U175 ( .A(n87), .B(N4961), .Z(n80) );
  CNR2IX1 U176 ( .B(N115), .A(N114), .Z(n87) );
  CAOR2X1 U177 ( .A(write_ptr[4]), .B(N213), .C(N218), .D(n100), .Z(N2526) );
  CAOR2X1 U178 ( .A(write_ptr[3]), .B(N213), .C(N217), .D(n100), .Z(N2524) );
  CAOR2X1 U179 ( .A(write_ptr[2]), .B(N213), .C(N216), .D(n100), .Z(N2523) );
  CAOR2X1 U180 ( .A(write_ptr[1]), .B(N213), .C(N215), .D(n100), .Z(N2522) );
  CAOR2X1 U181 ( .A(write_ptr[0]), .B(N213), .C(N214), .D(n100), .Z(N2521) );
  CNR2X1 U185 ( .A(n84), .B(N210), .Z(N213) );
  CIVX1 U186 ( .A(n90), .Z(n84) );
  CNR2X1 U187 ( .A(N114), .B(N115), .Z(n90) );
  CAN2X1 U188 ( .A(out[61]), .B(N122), .Z(N209) );
  CAN2X1 U189 ( .A(out[60]), .B(N122), .Z(N208) );
  CAN2X1 U190 ( .A(out[59]), .B(N122), .Z(N207) );
  CAN2X1 U191 ( .A(out[58]), .B(N122), .Z(N206) );
  CAN2X1 U192 ( .A(out[57]), .B(N122), .Z(N205) );
  CAN2X1 U193 ( .A(out[56]), .B(N122), .Z(N204) );
  CAN2X1 U194 ( .A(out[55]), .B(N122), .Z(N203) );
  CAN2X1 U195 ( .A(out[54]), .B(N122), .Z(N202) );
  CAN2X1 U196 ( .A(out[53]), .B(N122), .Z(N201) );
  CAN2X1 U197 ( .A(out[52]), .B(N122), .Z(N200) );
  CAN2X1 U198 ( .A(out[51]), .B(N122), .Z(N199) );
  CAN2X1 U199 ( .A(out[50]), .B(N122), .Z(N198) );
  CAN2X1 U200 ( .A(out[49]), .B(N122), .Z(N197) );
  CAN2X1 U201 ( .A(out[48]), .B(N122), .Z(N196) );
  CAN2X1 U202 ( .A(out[47]), .B(N122), .Z(N195) );
  CAN2X1 U203 ( .A(out[46]), .B(N122), .Z(N194) );
  CAN2X1 U204 ( .A(out[45]), .B(N122), .Z(N193) );
  CAN2X1 U205 ( .A(out[44]), .B(N122), .Z(N192) );
  CAN2X1 U206 ( .A(out[43]), .B(N122), .Z(N191) );
  CAN2X1 U207 ( .A(out[42]), .B(N122), .Z(N190) );
  CAN2X1 U208 ( .A(out[41]), .B(N122), .Z(N189) );
  CAN2X1 U209 ( .A(out[40]), .B(N122), .Z(N188) );
  CAN2X1 U210 ( .A(out[39]), .B(N122), .Z(N187) );
  CAN2X1 U211 ( .A(out[38]), .B(N122), .Z(N186) );
  CAN2X1 U212 ( .A(out[37]), .B(N122), .Z(N185) );
  CAN2X1 U213 ( .A(out[36]), .B(N122), .Z(N184) );
  CAN2X1 U214 ( .A(out[35]), .B(N122), .Z(N183) );
  CAN2X1 U215 ( .A(out[34]), .B(N122), .Z(N182) );
  CAN2X1 U216 ( .A(out[33]), .B(N122), .Z(N181) );
  CAN2X1 U217 ( .A(out[32]), .B(N122), .Z(N180) );
  CAN2X1 U218 ( .A(out[31]), .B(N122), .Z(N179) );
  CAN2X1 U219 ( .A(out[30]), .B(N122), .Z(N178) );
  CAN2X1 U220 ( .A(out[29]), .B(N122), .Z(N177) );
  CAN2X1 U221 ( .A(out[28]), .B(N122), .Z(N176) );
  CAN2X1 U222 ( .A(out[27]), .B(N122), .Z(N175) );
  CAN2X1 U223 ( .A(out[26]), .B(N122), .Z(N174) );
  CAN2X1 U224 ( .A(out[25]), .B(N122), .Z(N173) );
  CAN2X1 U225 ( .A(out[24]), .B(N122), .Z(N172) );
  CAN2X1 U226 ( .A(out[23]), .B(N122), .Z(N171) );
  CAN2X1 U227 ( .A(out[22]), .B(N122), .Z(N170) );
  CAN2X1 U228 ( .A(out[21]), .B(N122), .Z(N169) );
  CAN2X1 U229 ( .A(out[20]), .B(N122), .Z(N168) );
  CAN2X1 U230 ( .A(out[19]), .B(N122), .Z(N167) );
  CAN2X1 U231 ( .A(out[18]), .B(N122), .Z(N166) );
  CAN2X1 U232 ( .A(out[17]), .B(N122), .Z(N165) );
  CAN2X1 U233 ( .A(out[16]), .B(N122), .Z(N164) );
  CAN2X1 U234 ( .A(out[15]), .B(N122), .Z(N163) );
  CAN2X1 U235 ( .A(out[14]), .B(N122), .Z(N162) );
  CAN2X1 U236 ( .A(out[13]), .B(N122), .Z(N161) );
  CAN2X1 U237 ( .A(out[12]), .B(N122), .Z(N160) );
  CAN2X1 U238 ( .A(out[11]), .B(N122), .Z(N159) );
  CAN2X1 U239 ( .A(out[10]), .B(N122), .Z(N158) );
  CAN2X1 U240 ( .A(out[9]), .B(N122), .Z(N157) );
  CAN2X1 U241 ( .A(out[8]), .B(N122), .Z(N156) );
  CAN2X1 U242 ( .A(out[7]), .B(N122), .Z(N155) );
  CAN2X1 U243 ( .A(out[6]), .B(N122), .Z(N154) );
  CAN2X1 U244 ( .A(out[5]), .B(N122), .Z(N153) );
  CAN2X1 U245 ( .A(out[4]), .B(N122), .Z(N152) );
  CAN2X1 U246 ( .A(out[3]), .B(N122), .Z(N151) );
  CAN2X1 U247 ( .A(out[2]), .B(N122), .Z(N150) );
  CAN2X1 U248 ( .A(out[1]), .B(N122), .Z(N149) );
  CAN2X1 U249 ( .A(out[0]), .B(N122), .Z(N148) );
  CAN2X1 U250 ( .A(datain), .B(N122), .Z(N147) );
  CAN2X1 U251 ( .A(N132), .B(N122), .Z(N146) );
  CAN2X1 U252 ( .A(N131), .B(N122), .Z(N145) );
  CAN2X1 U253 ( .A(N130), .B(N122), .Z(N144) );
  CAN2X1 U254 ( .A(N129), .B(N122), .Z(N143) );
  CAN2X1 U255 ( .A(N128), .B(N122), .Z(N142) );
  CAN2X1 U256 ( .A(N127), .B(N122), .Z(N141) );
  CAN2X1 U257 ( .A(N126), .B(N122), .Z(N140) );
  CND2X1 U258 ( .A(lastin), .B(n78), .Z(N124) );
  CND2X1 U259 ( .A(pushin), .B(n79), .Z(N121) );
  CMX2X1 U260 ( .A0(n2598), .A1(N147), .S(N5105), .Z(n2529) );
  CMX2X1 U261 ( .A0(n2597), .A1(N148), .S(N5105), .Z(n2528) );
  CMX2X1 U262 ( .A0(n2596), .A1(N149), .S(N5105), .Z(n2527) );
  CMX2X1 U263 ( .A0(n2595), .A1(N150), .S(N5105), .Z(n2526) );
  CMX2X1 U264 ( .A0(n2594), .A1(N151), .S(N5105), .Z(n2525) );
  CMX2X1 U265 ( .A0(n2593), .A1(N152), .S(N5105), .Z(n2524) );
  CMX2X1 U266 ( .A0(n2592), .A1(N153), .S(N5105), .Z(n2523) );
  CMX2X1 U267 ( .A0(n2591), .A1(N154), .S(N5105), .Z(n2522) );
  CMX2X1 U268 ( .A0(n2590), .A1(N155), .S(N5105), .Z(n2521) );
  CMX2X1 U269 ( .A0(n2589), .A1(N156), .S(N5105), .Z(n2520) );
  CMX2X1 U270 ( .A0(n2588), .A1(N157), .S(N5105), .Z(n2519) );
  CMX2X1 U271 ( .A0(n2587), .A1(N158), .S(N5105), .Z(n2518) );
  CMX2X1 U272 ( .A0(n2586), .A1(N159), .S(N5105), .Z(n2517) );
  CMX2X1 U273 ( .A0(n2585), .A1(N160), .S(N5105), .Z(n2516) );
  CMX2X1 U274 ( .A0(n2584), .A1(N161), .S(N5105), .Z(n2515) );
  CMX2X1 U275 ( .A0(n2583), .A1(N162), .S(N5105), .Z(n2514) );
  CMX2X1 U276 ( .A0(n2582), .A1(N163), .S(N5105), .Z(n2513) );
  CMX2X1 U277 ( .A0(n2581), .A1(N164), .S(N5105), .Z(n2512) );
  CMX2X1 U278 ( .A0(n2580), .A1(N165), .S(N5105), .Z(n2511) );
  CMX2X1 U279 ( .A0(n2579), .A1(N166), .S(N5105), .Z(n2510) );
  CMX2X1 U280 ( .A0(n2578), .A1(N167), .S(N5105), .Z(n2509) );
  CMX2X1 U281 ( .A0(n2577), .A1(N168), .S(N5105), .Z(n2508) );
  CMX2X1 U282 ( .A0(n2576), .A1(N169), .S(N5105), .Z(n2507) );
  CMX2X1 U283 ( .A0(n2575), .A1(N170), .S(N5105), .Z(n2506) );
  CMX2X1 U284 ( .A0(n2574), .A1(N171), .S(N5105), .Z(n2505) );
  CMX2X1 U285 ( .A0(n2573), .A1(N172), .S(N5105), .Z(n2504) );
  CMX2X1 U286 ( .A0(n2572), .A1(N173), .S(N5105), .Z(n2503) );
  CMX2X1 U287 ( .A0(n2571), .A1(N174), .S(N5105), .Z(n2502) );
  CMX2X1 U288 ( .A0(n2570), .A1(N175), .S(N5105), .Z(n2501) );
  CMX2X1 U289 ( .A0(n2569), .A1(N176), .S(N5105), .Z(n2500) );
  CMX2X1 U290 ( .A0(n2568), .A1(N177), .S(N5105), .Z(n2499) );
  CMX2X1 U291 ( .A0(n2567), .A1(N178), .S(N5105), .Z(n2498) );
  CMX2X1 U292 ( .A0(n2566), .A1(N179), .S(N5105), .Z(n2497) );
  CMX2X1 U293 ( .A0(n2565), .A1(N180), .S(N5105), .Z(n2496) );
  CMX2X1 U294 ( .A0(n2564), .A1(N181), .S(N5105), .Z(n2495) );
  CMX2X1 U295 ( .A0(n2563), .A1(N182), .S(N5105), .Z(n2494) );
  CMX2X1 U296 ( .A0(n2562), .A1(N183), .S(N5105), .Z(n2493) );
  CMX2X1 U297 ( .A0(n2561), .A1(N184), .S(N5105), .Z(n2492) );
  CMX2X1 U298 ( .A0(n2560), .A1(N185), .S(N5105), .Z(n2491) );
  CMX2X1 U299 ( .A0(n2559), .A1(N186), .S(N5105), .Z(n2490) );
  CMX2X1 U300 ( .A0(n2558), .A1(N187), .S(N5105), .Z(n2489) );
  CMX2X1 U301 ( .A0(n2557), .A1(N188), .S(N5105), .Z(n2488) );
  CMX2X1 U302 ( .A0(n2556), .A1(N189), .S(N5105), .Z(n2487) );
  CMX2X1 U303 ( .A0(n2555), .A1(N190), .S(N5105), .Z(n2486) );
  CMX2X1 U304 ( .A0(n2554), .A1(N191), .S(N5105), .Z(n2485) );
  CMX2X1 U305 ( .A0(n2553), .A1(N192), .S(N5105), .Z(n2484) );
  CMX2X1 U306 ( .A0(n2552), .A1(N193), .S(N5105), .Z(n2483) );
  CMX2X1 U307 ( .A0(n2551), .A1(N194), .S(N5105), .Z(n2482) );
  CMX2X1 U308 ( .A0(n2550), .A1(N195), .S(N5105), .Z(n2481) );
  CMX2X1 U309 ( .A0(n2549), .A1(N196), .S(N5105), .Z(n2480) );
  CMX2X1 U310 ( .A0(n2548), .A1(N197), .S(N5105), .Z(n2479) );
  CMX2X1 U311 ( .A0(n2547), .A1(N198), .S(N5105), .Z(n2478) );
  CMX2X1 U312 ( .A0(n2546), .A1(N199), .S(N5105), .Z(n2477) );
  CMX2X1 U313 ( .A0(n2545), .A1(N200), .S(N5105), .Z(n2476) );
  CMX2X1 U314 ( .A0(n2544), .A1(N201), .S(N5105), .Z(n2475) );
  CMX2X1 U315 ( .A0(n2543), .A1(N202), .S(N5105), .Z(n2474) );
  CMX2X1 U316 ( .A0(n2542), .A1(N203), .S(N5105), .Z(n2473) );
  CMX2X1 U317 ( .A0(n2541), .A1(N204), .S(N5105), .Z(n2472) );
  CMX2X1 U318 ( .A0(n2540), .A1(N205), .S(N5105), .Z(n2471) );
  CMX2X1 U319 ( .A0(n2539), .A1(N206), .S(N5105), .Z(n2470) );
  CMX2X1 U320 ( .A0(n2538), .A1(N207), .S(N5105), .Z(n2469) );
  CMX2X1 U321 ( .A0(n2537), .A1(N208), .S(N5105), .Z(n2468) );
  CMX2X1 U322 ( .A0(n2536), .A1(N209), .S(N5105), .Z(n2467) );
  CMX2X1 U323 ( .A0(n2599), .A1(N140), .S(N5105), .Z(n2466) );
  CMX2X1 U324 ( .A0(lout[1]), .A1(N141), .S(N5105), .Z(n2465) );
  CMX2X1 U325 ( .A0(lout[2]), .A1(N142), .S(N5105), .Z(n2464) );
  CMX2X1 U326 ( .A0(lout[3]), .A1(N143), .S(N5105), .Z(n2463) );
  CMX2X1 U327 ( .A0(lout[4]), .A1(N144), .S(N5105), .Z(n2462) );
  CMX2X1 U328 ( .A0(lout[5]), .A1(N145), .S(N5105), .Z(n2461) );
  CMX2X1 U329 ( .A0(lout[6]), .A1(N146), .S(N5105), .Z(n2460) );
  CMX2X1 U330 ( .A0(counter[0]), .A1(N2533), .S(N4961), .Z(n2459) );
  CMX2X1 U407 ( .A0(n2636), .A1(N2527), .S(N2531), .Z(n2382) );
  CMX2X1 U408 ( .A0(n2624), .A1(N2528), .S(N2531), .Z(n2381) );
  CMX2X1 U409 ( .A0(n2612), .A1(N2529), .S(N2531), .Z(n2380) );
  CMX2X1 U410 ( .A0(N41), .A1(N2530), .S(N2531), .Z(n2379) );
  CMX2X1 U411 ( .A0(N42), .A1(N2532), .S(N2531), .Z(n2378) );
  CMX2X1 U412 ( .A0(write_ptr[0]), .A1(N2521), .S(N2525), .Z(n2377) );
  CMX2X1 U413 ( .A0(write_ptr[1]), .A1(N2522), .S(N2525), .Z(n2376) );
  CMX2X1 U414 ( .A0(write_ptr[2]), .A1(N2523), .S(N2525), .Z(n2375) );
  CMX2X1 U415 ( .A0(write_ptr[3]), .A1(N2524), .S(N2525), .Z(n2374) );
  CMX2X1 U416 ( .A0(write_ptr[4]), .A1(N2526), .S(N2525), .Z(n2373) );
  serial_DW01_inc_3 r182 ( .A({lout[6:1], n2599}), .SUM({N132, N131, N130, 
        N129, N128, N127, N126}) );
  CHA1X1 \add_116/U1_1_1  ( .A(counter[1]), .B(counter[0]), .CO(
        \add_116/carry[2] ), .S(N231) );
  CHA1X1 \add_116/U1_1_2  ( .A(counter[2]), .B(\add_116/carry[2] ), .CO(
        \add_116/carry[3] ), .S(N232) );
  CHA1X1 \add_116/U1_1_3  ( .A(counter[3]), .B(\add_116/carry[3] ), .CO(
        \add_116/carry[4] ), .S(N233) );
  CHA1X1 \r184/U1_1_1  ( .A(n2624), .B(n2636), .CO(\r184/carry[2] ), .S(N220)
         );
  CHA1X1 \r184/U1_1_2  ( .A(n2612), .B(\r184/carry[2] ), .CO(\r184/carry[3] ), 
        .S(N221) );
  CHA1X1 \r184/U1_1_3  ( .A(N41), .B(\r184/carry[3] ), .CO(\r184/carry[4] ), 
        .S(N222) );
  CHA1X1 \r183/U1_1_1  ( .A(write_ptr[1]), .B(write_ptr[0]), .CO(
        \r183/carry[2] ), .S(N215) );
  CHA1X1 \r183/U1_1_2  ( .A(write_ptr[2]), .B(\r183/carry[2] ), .CO(
        \r183/carry[3] ), .S(N216) );
  CHA1X1 \r183/U1_1_3  ( .A(write_ptr[3]), .B(\r183/carry[3] ), .CO(
        \r183/carry[4] ), .S(N217) );
  CHA1XL \add_116/U1_1_4  ( .A(counter[4]), .B(\add_116/carry[4] ), .CO(
        \add_116/carry[5] ), .S(N234) );
  CIVX1 \stopout_reg/U7  ( .A(pullout), .Z(n2609) );
  CFD4QXL stopout_reg ( .D(n2608), .CP(clk), .SD(n77), .Q(stopout) );
  CIVX1 \read_reg/U5  ( .A(stopout), .Z(n2607) );
  CFD2QXL read_reg ( .D(n2606), .CP(clk), .CD(n77), .Q(read) );
  CFD2QXL write_reg ( .D(N123), .CP(clk), .CD(n77), .Q(write) );
  CFD1QXL \memory_reg[31][70]  ( .D(n101), .CP(clk), .Q(\memory[31][70] ) );
  CFD1QXL \memory_reg[31][69]  ( .D(n102), .CP(clk), .Q(\memory[31][69] ) );
  CFD1QXL \memory_reg[31][68]  ( .D(n103), .CP(clk), .Q(\memory[31][68] ) );
  CFD1QXL \memory_reg[31][67]  ( .D(n104), .CP(clk), .Q(\memory[31][67] ) );
  CFD1QXL \memory_reg[31][66]  ( .D(n105), .CP(clk), .Q(\memory[31][66] ) );
  CFD1QXL \memory_reg[31][65]  ( .D(n106), .CP(clk), .Q(\memory[31][65] ) );
  CFD1QXL \memory_reg[31][64]  ( .D(n107), .CP(clk), .Q(\memory[31][64] ) );
  CFD1QXL \memory_reg[30][70]  ( .D(n172), .CP(clk), .Q(\memory[30][70] ) );
  CFD1QXL \memory_reg[30][69]  ( .D(n173), .CP(clk), .Q(\memory[30][69] ) );
  CFD1QXL \memory_reg[30][68]  ( .D(n174), .CP(clk), .Q(\memory[30][68] ) );
  CFD1QXL \memory_reg[30][67]  ( .D(n175), .CP(clk), .Q(\memory[30][67] ) );
  CFD1QXL \memory_reg[30][66]  ( .D(n176), .CP(clk), .Q(\memory[30][66] ) );
  CFD1QXL \memory_reg[30][65]  ( .D(n177), .CP(clk), .Q(\memory[30][65] ) );
  CFD1QXL \memory_reg[30][64]  ( .D(n178), .CP(clk), .Q(\memory[30][64] ) );
  CFD1QXL \memory_reg[29][70]  ( .D(n243), .CP(clk), .Q(\memory[29][70] ) );
  CFD1QXL \memory_reg[29][69]  ( .D(n244), .CP(clk), .Q(\memory[29][69] ) );
  CFD1QXL \memory_reg[29][68]  ( .D(n245), .CP(clk), .Q(\memory[29][68] ) );
  CFD1QXL \memory_reg[29][67]  ( .D(n246), .CP(clk), .Q(\memory[29][67] ) );
  CFD1QXL \memory_reg[29][66]  ( .D(n247), .CP(clk), .Q(\memory[29][66] ) );
  CFD1QXL \memory_reg[29][65]  ( .D(n248), .CP(clk), .Q(\memory[29][65] ) );
  CFD1QXL \memory_reg[29][64]  ( .D(n249), .CP(clk), .Q(\memory[29][64] ) );
  CFD1QXL \memory_reg[28][70]  ( .D(n314), .CP(clk), .Q(\memory[28][70] ) );
  CFD1QXL \memory_reg[28][69]  ( .D(n315), .CP(clk), .Q(\memory[28][69] ) );
  CFD1QXL \memory_reg[28][68]  ( .D(n316), .CP(clk), .Q(\memory[28][68] ) );
  CFD1QXL \memory_reg[28][67]  ( .D(n317), .CP(clk), .Q(\memory[28][67] ) );
  CFD1QXL \memory_reg[28][66]  ( .D(n318), .CP(clk), .Q(\memory[28][66] ) );
  CFD1QXL \memory_reg[28][65]  ( .D(n319), .CP(clk), .Q(\memory[28][65] ) );
  CFD1QXL \memory_reg[28][64]  ( .D(n320), .CP(clk), .Q(\memory[28][64] ) );
  CFD1QXL \memory_reg[27][70]  ( .D(n385), .CP(clk), .Q(\memory[27][70] ) );
  CFD1QXL \memory_reg[27][69]  ( .D(n386), .CP(clk), .Q(\memory[27][69] ) );
  CFD1QXL \memory_reg[27][68]  ( .D(n387), .CP(clk), .Q(\memory[27][68] ) );
  CFD1QXL \memory_reg[27][67]  ( .D(n388), .CP(clk), .Q(\memory[27][67] ) );
  CFD1QXL \memory_reg[27][66]  ( .D(n389), .CP(clk), .Q(\memory[27][66] ) );
  CFD1QXL \memory_reg[27][65]  ( .D(n390), .CP(clk), .Q(\memory[27][65] ) );
  CFD1QXL \memory_reg[27][64]  ( .D(n391), .CP(clk), .Q(\memory[27][64] ) );
  CFD1QXL \memory_reg[26][70]  ( .D(n456), .CP(clk), .Q(\memory[26][70] ) );
  CFD1QXL \memory_reg[26][69]  ( .D(n457), .CP(clk), .Q(\memory[26][69] ) );
  CFD1QXL \memory_reg[26][68]  ( .D(n458), .CP(clk), .Q(\memory[26][68] ) );
  CFD1QXL \memory_reg[26][67]  ( .D(n459), .CP(clk), .Q(\memory[26][67] ) );
  CFD1QXL \memory_reg[26][66]  ( .D(n460), .CP(clk), .Q(\memory[26][66] ) );
  CFD1QXL \memory_reg[26][65]  ( .D(n461), .CP(clk), .Q(\memory[26][65] ) );
  CFD1QXL \memory_reg[26][64]  ( .D(n462), .CP(clk), .Q(\memory[26][64] ) );
  CFD1QXL \memory_reg[25][70]  ( .D(n527), .CP(clk), .Q(\memory[25][70] ) );
  CFD1QXL \memory_reg[25][69]  ( .D(n528), .CP(clk), .Q(\memory[25][69] ) );
  CFD1QXL \memory_reg[25][68]  ( .D(n529), .CP(clk), .Q(\memory[25][68] ) );
  CFD1QXL \memory_reg[25][67]  ( .D(n530), .CP(clk), .Q(\memory[25][67] ) );
  CFD1QXL \memory_reg[25][66]  ( .D(n531), .CP(clk), .Q(\memory[25][66] ) );
  CFD1QXL \memory_reg[25][65]  ( .D(n532), .CP(clk), .Q(\memory[25][65] ) );
  CFD1QXL \memory_reg[25][64]  ( .D(n533), .CP(clk), .Q(\memory[25][64] ) );
  CFD1QXL \memory_reg[24][70]  ( .D(n598), .CP(clk), .Q(\memory[24][70] ) );
  CFD1QXL \memory_reg[24][69]  ( .D(n599), .CP(clk), .Q(\memory[24][69] ) );
  CFD1QXL \memory_reg[24][68]  ( .D(n600), .CP(clk), .Q(\memory[24][68] ) );
  CFD1QXL \memory_reg[24][67]  ( .D(n601), .CP(clk), .Q(\memory[24][67] ) );
  CFD1QXL \memory_reg[24][66]  ( .D(n602), .CP(clk), .Q(\memory[24][66] ) );
  CFD1QXL \memory_reg[24][65]  ( .D(n603), .CP(clk), .Q(\memory[24][65] ) );
  CFD1QXL \memory_reg[24][64]  ( .D(n604), .CP(clk), .Q(\memory[24][64] ) );
  CFD1QXL \memory_reg[23][70]  ( .D(n669), .CP(clk), .Q(\memory[23][70] ) );
  CFD1QXL \memory_reg[23][69]  ( .D(n670), .CP(clk), .Q(\memory[23][69] ) );
  CFD1QXL \memory_reg[23][68]  ( .D(n671), .CP(clk), .Q(\memory[23][68] ) );
  CFD1QXL \memory_reg[23][67]  ( .D(n672), .CP(clk), .Q(\memory[23][67] ) );
  CFD1QXL \memory_reg[23][66]  ( .D(n673), .CP(clk), .Q(\memory[23][66] ) );
  CFD1QXL \memory_reg[23][65]  ( .D(n674), .CP(clk), .Q(\memory[23][65] ) );
  CFD1QXL \memory_reg[23][64]  ( .D(n675), .CP(clk), .Q(\memory[23][64] ) );
  CFD1QXL \memory_reg[22][70]  ( .D(n740), .CP(clk), .Q(\memory[22][70] ) );
  CFD1QXL \memory_reg[22][69]  ( .D(n741), .CP(clk), .Q(\memory[22][69] ) );
  CFD1QXL \memory_reg[22][68]  ( .D(n742), .CP(clk), .Q(\memory[22][68] ) );
  CFD1QXL \memory_reg[22][67]  ( .D(n743), .CP(clk), .Q(\memory[22][67] ) );
  CFD1QXL \memory_reg[22][66]  ( .D(n744), .CP(clk), .Q(\memory[22][66] ) );
  CFD1QXL \memory_reg[22][65]  ( .D(n745), .CP(clk), .Q(\memory[22][65] ) );
  CFD1QXL \memory_reg[22][64]  ( .D(n746), .CP(clk), .Q(\memory[22][64] ) );
  CFD1QXL \memory_reg[21][70]  ( .D(n811), .CP(clk), .Q(\memory[21][70] ) );
  CFD1QXL \memory_reg[21][69]  ( .D(n812), .CP(clk), .Q(\memory[21][69] ) );
  CFD1QXL \memory_reg[21][68]  ( .D(n813), .CP(clk), .Q(\memory[21][68] ) );
  CFD1QXL \memory_reg[21][67]  ( .D(n814), .CP(clk), .Q(\memory[21][67] ) );
  CFD1QXL \memory_reg[21][66]  ( .D(n815), .CP(clk), .Q(\memory[21][66] ) );
  CFD1QXL \memory_reg[21][65]  ( .D(n816), .CP(clk), .Q(\memory[21][65] ) );
  CFD1QXL \memory_reg[21][64]  ( .D(n817), .CP(clk), .Q(\memory[21][64] ) );
  CFD1QXL \memory_reg[20][70]  ( .D(n882), .CP(clk), .Q(\memory[20][70] ) );
  CFD1QXL \memory_reg[20][69]  ( .D(n883), .CP(clk), .Q(\memory[20][69] ) );
  CFD1QXL \memory_reg[20][68]  ( .D(n884), .CP(clk), .Q(\memory[20][68] ) );
  CFD1QXL \memory_reg[20][67]  ( .D(n885), .CP(clk), .Q(\memory[20][67] ) );
  CFD1QXL \memory_reg[20][66]  ( .D(n886), .CP(clk), .Q(\memory[20][66] ) );
  CFD1QXL \memory_reg[20][65]  ( .D(n887), .CP(clk), .Q(\memory[20][65] ) );
  CFD1QXL \memory_reg[20][64]  ( .D(n888), .CP(clk), .Q(\memory[20][64] ) );
  CFD1QXL \memory_reg[19][70]  ( .D(n953), .CP(clk), .Q(\memory[19][70] ) );
  CFD1QXL \memory_reg[19][69]  ( .D(n954), .CP(clk), .Q(\memory[19][69] ) );
  CFD1QXL \memory_reg[19][68]  ( .D(n955), .CP(clk), .Q(\memory[19][68] ) );
  CFD1QXL \memory_reg[19][67]  ( .D(n956), .CP(clk), .Q(\memory[19][67] ) );
  CFD1QXL \memory_reg[19][66]  ( .D(n957), .CP(clk), .Q(\memory[19][66] ) );
  CFD1QXL \memory_reg[19][65]  ( .D(n958), .CP(clk), .Q(\memory[19][65] ) );
  CFD1QXL \memory_reg[19][64]  ( .D(n959), .CP(clk), .Q(\memory[19][64] ) );
  CFD1QXL \memory_reg[18][70]  ( .D(n1024), .CP(clk), .Q(\memory[18][70] ) );
  CFD1QXL \memory_reg[18][69]  ( .D(n1025), .CP(clk), .Q(\memory[18][69] ) );
  CFD1QXL \memory_reg[18][68]  ( .D(n1026), .CP(clk), .Q(\memory[18][68] ) );
  CFD1QXL \memory_reg[18][67]  ( .D(n1027), .CP(clk), .Q(\memory[18][67] ) );
  CFD1QXL \memory_reg[18][66]  ( .D(n1028), .CP(clk), .Q(\memory[18][66] ) );
  CFD1QXL \memory_reg[18][65]  ( .D(n1029), .CP(clk), .Q(\memory[18][65] ) );
  CFD1QXL \memory_reg[18][64]  ( .D(n1030), .CP(clk), .Q(\memory[18][64] ) );
  CFD1QXL \memory_reg[17][70]  ( .D(n1095), .CP(clk), .Q(\memory[17][70] ) );
  CFD1QXL \memory_reg[17][69]  ( .D(n1096), .CP(clk), .Q(\memory[17][69] ) );
  CFD1QXL \memory_reg[17][68]  ( .D(n1097), .CP(clk), .Q(\memory[17][68] ) );
  CFD1QXL \memory_reg[17][67]  ( .D(n1098), .CP(clk), .Q(\memory[17][67] ) );
  CFD1QXL \memory_reg[17][66]  ( .D(n1099), .CP(clk), .Q(\memory[17][66] ) );
  CFD1QXL \memory_reg[17][65]  ( .D(n1100), .CP(clk), .Q(\memory[17][65] ) );
  CFD1QXL \memory_reg[17][64]  ( .D(n1101), .CP(clk), .Q(\memory[17][64] ) );
  CFD1QXL \memory_reg[16][70]  ( .D(n1166), .CP(clk), .Q(\memory[16][70] ) );
  CFD1QXL \memory_reg[16][69]  ( .D(n1167), .CP(clk), .Q(\memory[16][69] ) );
  CFD1QXL \memory_reg[16][68]  ( .D(n1168), .CP(clk), .Q(\memory[16][68] ) );
  CFD1QXL \memory_reg[16][67]  ( .D(n1169), .CP(clk), .Q(\memory[16][67] ) );
  CFD1QXL \memory_reg[16][66]  ( .D(n1170), .CP(clk), .Q(\memory[16][66] ) );
  CFD1QXL \memory_reg[16][65]  ( .D(n1171), .CP(clk), .Q(\memory[16][65] ) );
  CFD1QXL \memory_reg[16][64]  ( .D(n1172), .CP(clk), .Q(\memory[16][64] ) );
  CFD1QXL \memory_reg[15][70]  ( .D(n1237), .CP(clk), .Q(\memory[15][70] ) );
  CFD1QXL \memory_reg[15][69]  ( .D(n1238), .CP(clk), .Q(\memory[15][69] ) );
  CFD1QXL \memory_reg[15][68]  ( .D(n1239), .CP(clk), .Q(\memory[15][68] ) );
  CFD1QXL \memory_reg[15][67]  ( .D(n1240), .CP(clk), .Q(\memory[15][67] ) );
  CFD1QXL \memory_reg[15][66]  ( .D(n1241), .CP(clk), .Q(\memory[15][66] ) );
  CFD1QXL \memory_reg[15][65]  ( .D(n1242), .CP(clk), .Q(\memory[15][65] ) );
  CFD1QXL \memory_reg[15][64]  ( .D(n1243), .CP(clk), .Q(\memory[15][64] ) );
  CFD1QXL \memory_reg[14][70]  ( .D(n1308), .CP(clk), .Q(\memory[14][70] ) );
  CFD1QXL \memory_reg[14][69]  ( .D(n1309), .CP(clk), .Q(\memory[14][69] ) );
  CFD1QXL \memory_reg[14][68]  ( .D(n1310), .CP(clk), .Q(\memory[14][68] ) );
  CFD1QXL \memory_reg[14][67]  ( .D(n1311), .CP(clk), .Q(\memory[14][67] ) );
  CFD1QXL \memory_reg[14][66]  ( .D(n1312), .CP(clk), .Q(\memory[14][66] ) );
  CFD1QXL \memory_reg[14][65]  ( .D(n1313), .CP(clk), .Q(\memory[14][65] ) );
  CFD1QXL \memory_reg[14][64]  ( .D(n1314), .CP(clk), .Q(\memory[14][64] ) );
  CFD1QXL \memory_reg[13][70]  ( .D(n1379), .CP(clk), .Q(\memory[13][70] ) );
  CFD1QXL \memory_reg[13][69]  ( .D(n1380), .CP(clk), .Q(\memory[13][69] ) );
  CFD1QXL \memory_reg[13][68]  ( .D(n1381), .CP(clk), .Q(\memory[13][68] ) );
  CFD1QXL \memory_reg[13][67]  ( .D(n1382), .CP(clk), .Q(\memory[13][67] ) );
  CFD1QXL \memory_reg[13][66]  ( .D(n1383), .CP(clk), .Q(\memory[13][66] ) );
  CFD1QXL \memory_reg[13][65]  ( .D(n1384), .CP(clk), .Q(\memory[13][65] ) );
  CFD1QXL \memory_reg[13][64]  ( .D(n1385), .CP(clk), .Q(\memory[13][64] ) );
  CFD1QXL \memory_reg[12][70]  ( .D(n1450), .CP(clk), .Q(\memory[12][70] ) );
  CFD1QXL \memory_reg[12][69]  ( .D(n1451), .CP(clk), .Q(\memory[12][69] ) );
  CFD1QXL \memory_reg[12][68]  ( .D(n1452), .CP(clk), .Q(\memory[12][68] ) );
  CFD1QXL \memory_reg[12][67]  ( .D(n1453), .CP(clk), .Q(\memory[12][67] ) );
  CFD1QXL \memory_reg[12][66]  ( .D(n1454), .CP(clk), .Q(\memory[12][66] ) );
  CFD1QXL \memory_reg[12][65]  ( .D(n1455), .CP(clk), .Q(\memory[12][65] ) );
  CFD1QXL \memory_reg[12][64]  ( .D(n1456), .CP(clk), .Q(\memory[12][64] ) );
  CFD1QXL \memory_reg[11][70]  ( .D(n1521), .CP(clk), .Q(\memory[11][70] ) );
  CFD1QXL \memory_reg[11][69]  ( .D(n1522), .CP(clk), .Q(\memory[11][69] ) );
  CFD1QXL \memory_reg[11][68]  ( .D(n1523), .CP(clk), .Q(\memory[11][68] ) );
  CFD1QXL \memory_reg[11][67]  ( .D(n1524), .CP(clk), .Q(\memory[11][67] ) );
  CFD1QXL \memory_reg[11][66]  ( .D(n1525), .CP(clk), .Q(\memory[11][66] ) );
  CFD1QXL \memory_reg[11][65]  ( .D(n1526), .CP(clk), .Q(\memory[11][65] ) );
  CFD1QXL \memory_reg[11][64]  ( .D(n1527), .CP(clk), .Q(\memory[11][64] ) );
  CFD1QXL \memory_reg[10][70]  ( .D(n1592), .CP(clk), .Q(\memory[10][70] ) );
  CFD1QXL \memory_reg[10][69]  ( .D(n1593), .CP(clk), .Q(\memory[10][69] ) );
  CFD1QXL \memory_reg[10][68]  ( .D(n1594), .CP(clk), .Q(\memory[10][68] ) );
  CFD1QXL \memory_reg[10][67]  ( .D(n1595), .CP(clk), .Q(\memory[10][67] ) );
  CFD1QXL \memory_reg[10][66]  ( .D(n1596), .CP(clk), .Q(\memory[10][66] ) );
  CFD1QXL \memory_reg[10][65]  ( .D(n1597), .CP(clk), .Q(\memory[10][65] ) );
  CFD1QXL \memory_reg[10][64]  ( .D(n1598), .CP(clk), .Q(\memory[10][64] ) );
  CFD1QXL \memory_reg[9][70]  ( .D(n1663), .CP(clk), .Q(\memory[9][70] ) );
  CFD1QXL \memory_reg[9][69]  ( .D(n1664), .CP(clk), .Q(\memory[9][69] ) );
  CFD1QXL \memory_reg[9][68]  ( .D(n1665), .CP(clk), .Q(\memory[9][68] ) );
  CFD1QXL \memory_reg[9][67]  ( .D(n1666), .CP(clk), .Q(\memory[9][67] ) );
  CFD1QXL \memory_reg[9][66]  ( .D(n1667), .CP(clk), .Q(\memory[9][66] ) );
  CFD1QXL \memory_reg[9][65]  ( .D(n1668), .CP(clk), .Q(\memory[9][65] ) );
  CFD1QXL \memory_reg[9][64]  ( .D(n1669), .CP(clk), .Q(\memory[9][64] ) );
  CFD1QXL \memory_reg[8][70]  ( .D(n1734), .CP(clk), .Q(\memory[8][70] ) );
  CFD1QXL \memory_reg[8][69]  ( .D(n1735), .CP(clk), .Q(\memory[8][69] ) );
  CFD1QXL \memory_reg[8][68]  ( .D(n1736), .CP(clk), .Q(\memory[8][68] ) );
  CFD1QXL \memory_reg[8][67]  ( .D(n1737), .CP(clk), .Q(\memory[8][67] ) );
  CFD1QXL \memory_reg[8][66]  ( .D(n1738), .CP(clk), .Q(\memory[8][66] ) );
  CFD1QXL \memory_reg[8][65]  ( .D(n1739), .CP(clk), .Q(\memory[8][65] ) );
  CFD1QXL \memory_reg[8][64]  ( .D(n1740), .CP(clk), .Q(\memory[8][64] ) );
  CFD1QXL \memory_reg[7][70]  ( .D(n1805), .CP(clk), .Q(\memory[7][70] ) );
  CFD1QXL \memory_reg[7][69]  ( .D(n1806), .CP(clk), .Q(\memory[7][69] ) );
  CFD1QXL \memory_reg[7][68]  ( .D(n1807), .CP(clk), .Q(\memory[7][68] ) );
  CFD1QXL \memory_reg[7][67]  ( .D(n1808), .CP(clk), .Q(\memory[7][67] ) );
  CFD1QXL \memory_reg[7][66]  ( .D(n1809), .CP(clk), .Q(\memory[7][66] ) );
  CFD1QXL \memory_reg[7][65]  ( .D(n1810), .CP(clk), .Q(\memory[7][65] ) );
  CFD1QXL \memory_reg[7][64]  ( .D(n1811), .CP(clk), .Q(\memory[7][64] ) );
  CFD1QXL \memory_reg[6][70]  ( .D(n1876), .CP(clk), .Q(\memory[6][70] ) );
  CFD1QXL \memory_reg[6][69]  ( .D(n1877), .CP(clk), .Q(\memory[6][69] ) );
  CFD1QXL \memory_reg[6][68]  ( .D(n1878), .CP(clk), .Q(\memory[6][68] ) );
  CFD1QXL \memory_reg[6][67]  ( .D(n1879), .CP(clk), .Q(\memory[6][67] ) );
  CFD1QXL \memory_reg[6][66]  ( .D(n1880), .CP(clk), .Q(\memory[6][66] ) );
  CFD1QXL \memory_reg[6][65]  ( .D(n1881), .CP(clk), .Q(\memory[6][65] ) );
  CFD1QXL \memory_reg[6][64]  ( .D(n1882), .CP(clk), .Q(\memory[6][64] ) );
  CFD1QXL \memory_reg[5][70]  ( .D(n1947), .CP(clk), .Q(\memory[5][70] ) );
  CFD1QXL \memory_reg[5][69]  ( .D(n1948), .CP(clk), .Q(\memory[5][69] ) );
  CFD1QXL \memory_reg[5][68]  ( .D(n1949), .CP(clk), .Q(\memory[5][68] ) );
  CFD1QXL \memory_reg[5][67]  ( .D(n1950), .CP(clk), .Q(\memory[5][67] ) );
  CFD1QXL \memory_reg[5][66]  ( .D(n1951), .CP(clk), .Q(\memory[5][66] ) );
  CFD1QXL \memory_reg[5][65]  ( .D(n1952), .CP(clk), .Q(\memory[5][65] ) );
  CFD1QXL \memory_reg[5][64]  ( .D(n1953), .CP(clk), .Q(\memory[5][64] ) );
  CFD1QXL \memory_reg[4][70]  ( .D(n2018), .CP(clk), .Q(\memory[4][70] ) );
  CFD1QXL \memory_reg[4][69]  ( .D(n2019), .CP(clk), .Q(\memory[4][69] ) );
  CFD1QXL \memory_reg[4][68]  ( .D(n2020), .CP(clk), .Q(\memory[4][68] ) );
  CFD1QXL \memory_reg[4][67]  ( .D(n2021), .CP(clk), .Q(\memory[4][67] ) );
  CFD1QXL \memory_reg[4][66]  ( .D(n2022), .CP(clk), .Q(\memory[4][66] ) );
  CFD1QXL \memory_reg[4][65]  ( .D(n2023), .CP(clk), .Q(\memory[4][65] ) );
  CFD1QXL \memory_reg[4][64]  ( .D(n2024), .CP(clk), .Q(\memory[4][64] ) );
  CFD1QXL \memory_reg[3][70]  ( .D(n2089), .CP(clk), .Q(\memory[3][70] ) );
  CFD1QXL \memory_reg[3][69]  ( .D(n2090), .CP(clk), .Q(\memory[3][69] ) );
  CFD1QXL \memory_reg[3][68]  ( .D(n2091), .CP(clk), .Q(\memory[3][68] ) );
  CFD1QXL \memory_reg[3][67]  ( .D(n2092), .CP(clk), .Q(\memory[3][67] ) );
  CFD1QXL \memory_reg[3][66]  ( .D(n2093), .CP(clk), .Q(\memory[3][66] ) );
  CFD1QXL \memory_reg[3][65]  ( .D(n2094), .CP(clk), .Q(\memory[3][65] ) );
  CFD1QXL \memory_reg[3][64]  ( .D(n2095), .CP(clk), .Q(\memory[3][64] ) );
  CFD1QXL \memory_reg[2][70]  ( .D(n2160), .CP(clk), .Q(\memory[2][70] ) );
  CFD1QXL \memory_reg[2][69]  ( .D(n2161), .CP(clk), .Q(\memory[2][69] ) );
  CFD1QXL \memory_reg[2][68]  ( .D(n2162), .CP(clk), .Q(\memory[2][68] ) );
  CFD1QXL \memory_reg[2][67]  ( .D(n2163), .CP(clk), .Q(\memory[2][67] ) );
  CFD1QXL \memory_reg[2][66]  ( .D(n2164), .CP(clk), .Q(\memory[2][66] ) );
  CFD1QXL \memory_reg[2][65]  ( .D(n2165), .CP(clk), .Q(\memory[2][65] ) );
  CFD1QXL \memory_reg[2][64]  ( .D(n2166), .CP(clk), .Q(\memory[2][64] ) );
  CFD1QXL \memory_reg[1][70]  ( .D(n2231), .CP(clk), .Q(\memory[1][70] ) );
  CFD1QXL \memory_reg[1][69]  ( .D(n2232), .CP(clk), .Q(\memory[1][69] ) );
  CFD1QXL \memory_reg[1][68]  ( .D(n2233), .CP(clk), .Q(\memory[1][68] ) );
  CFD1QXL \memory_reg[1][67]  ( .D(n2234), .CP(clk), .Q(\memory[1][67] ) );
  CFD1QXL \memory_reg[1][66]  ( .D(n2235), .CP(clk), .Q(\memory[1][66] ) );
  CFD1QXL \memory_reg[1][65]  ( .D(n2236), .CP(clk), .Q(\memory[1][65] ) );
  CFD1QXL \memory_reg[1][64]  ( .D(n2237), .CP(clk), .Q(\memory[1][64] ) );
  CFD1QXL \memory_reg[0][70]  ( .D(n2302), .CP(clk), .Q(\memory[0][70] ) );
  CFD1QXL \memory_reg[0][69]  ( .D(n2303), .CP(clk), .Q(\memory[0][69] ) );
  CFD1QXL \memory_reg[0][68]  ( .D(n2304), .CP(clk), .Q(\memory[0][68] ) );
  CFD1QXL \memory_reg[0][67]  ( .D(n2305), .CP(clk), .Q(\memory[0][67] ) );
  CFD1QXL \memory_reg[0][66]  ( .D(n2306), .CP(clk), .Q(\memory[0][66] ) );
  CFD1QXL \memory_reg[0][65]  ( .D(n2307), .CP(clk), .Q(\memory[0][65] ) );
  CFD1QXL \memory_reg[0][64]  ( .D(n2308), .CP(clk), .Q(\memory[0][64] ) );
  CFD1QXL \memory_reg[31][63]  ( .D(n108), .CP(clk), .Q(\memory[31][63] ) );
  CFD1QXL \memory_reg[31][62]  ( .D(n109), .CP(clk), .Q(\memory[31][62] ) );
  CFD1QXL \memory_reg[31][61]  ( .D(n110), .CP(clk), .Q(\memory[31][61] ) );
  CFD1QXL \memory_reg[31][60]  ( .D(n111), .CP(clk), .Q(\memory[31][60] ) );
  CFD1QXL \memory_reg[31][59]  ( .D(n112), .CP(clk), .Q(\memory[31][59] ) );
  CFD1QXL \memory_reg[31][58]  ( .D(n113), .CP(clk), .Q(\memory[31][58] ) );
  CFD1QXL \memory_reg[31][57]  ( .D(n114), .CP(clk), .Q(\memory[31][57] ) );
  CFD1QXL \memory_reg[31][56]  ( .D(n115), .CP(clk), .Q(\memory[31][56] ) );
  CFD1QXL \memory_reg[31][55]  ( .D(n116), .CP(clk), .Q(\memory[31][55] ) );
  CFD1QXL \memory_reg[31][54]  ( .D(n117), .CP(clk), .Q(\memory[31][54] ) );
  CFD1QXL \memory_reg[31][53]  ( .D(n118), .CP(clk), .Q(\memory[31][53] ) );
  CFD1QXL \memory_reg[31][52]  ( .D(n119), .CP(clk), .Q(\memory[31][52] ) );
  CFD1QXL \memory_reg[31][51]  ( .D(n120), .CP(clk), .Q(\memory[31][51] ) );
  CFD1QXL \memory_reg[31][50]  ( .D(n121), .CP(clk), .Q(\memory[31][50] ) );
  CFD1QXL \memory_reg[31][49]  ( .D(n122), .CP(clk), .Q(\memory[31][49] ) );
  CFD1QXL \memory_reg[31][48]  ( .D(n123), .CP(clk), .Q(\memory[31][48] ) );
  CFD1QXL \memory_reg[31][47]  ( .D(n124), .CP(clk), .Q(\memory[31][47] ) );
  CFD1QXL \memory_reg[31][46]  ( .D(n125), .CP(clk), .Q(\memory[31][46] ) );
  CFD1QXL \memory_reg[31][45]  ( .D(n126), .CP(clk), .Q(\memory[31][45] ) );
  CFD1QXL \memory_reg[31][44]  ( .D(n127), .CP(clk), .Q(\memory[31][44] ) );
  CFD1QXL \memory_reg[31][43]  ( .D(n128), .CP(clk), .Q(\memory[31][43] ) );
  CFD1QXL \memory_reg[31][42]  ( .D(n129), .CP(clk), .Q(\memory[31][42] ) );
  CFD1QXL \memory_reg[31][41]  ( .D(n130), .CP(clk), .Q(\memory[31][41] ) );
  CFD1QXL \memory_reg[31][40]  ( .D(n131), .CP(clk), .Q(\memory[31][40] ) );
  CFD1QXL \memory_reg[31][39]  ( .D(n132), .CP(clk), .Q(\memory[31][39] ) );
  CFD1QXL \memory_reg[31][38]  ( .D(n133), .CP(clk), .Q(\memory[31][38] ) );
  CFD1QXL \memory_reg[31][37]  ( .D(n134), .CP(clk), .Q(\memory[31][37] ) );
  CFD1QXL \memory_reg[31][36]  ( .D(n135), .CP(clk), .Q(\memory[31][36] ) );
  CFD1QXL \memory_reg[31][35]  ( .D(n136), .CP(clk), .Q(\memory[31][35] ) );
  CFD1QXL \memory_reg[31][34]  ( .D(n137), .CP(clk), .Q(\memory[31][34] ) );
  CFD1QXL \memory_reg[31][33]  ( .D(n138), .CP(clk), .Q(\memory[31][33] ) );
  CFD1QXL \memory_reg[31][32]  ( .D(n139), .CP(clk), .Q(\memory[31][32] ) );
  CFD1QXL \memory_reg[31][31]  ( .D(n140), .CP(clk), .Q(\memory[31][31] ) );
  CFD1QXL \memory_reg[31][30]  ( .D(n141), .CP(clk), .Q(\memory[31][30] ) );
  CFD1QXL \memory_reg[31][29]  ( .D(n142), .CP(clk), .Q(\memory[31][29] ) );
  CFD1QXL \memory_reg[31][28]  ( .D(n143), .CP(clk), .Q(\memory[31][28] ) );
  CFD1QXL \memory_reg[31][27]  ( .D(n144), .CP(clk), .Q(\memory[31][27] ) );
  CFD1QXL \memory_reg[31][26]  ( .D(n145), .CP(clk), .Q(\memory[31][26] ) );
  CFD1QXL \memory_reg[31][25]  ( .D(n146), .CP(clk), .Q(\memory[31][25] ) );
  CFD1QXL \memory_reg[31][24]  ( .D(n147), .CP(clk), .Q(\memory[31][24] ) );
  CFD1QXL \memory_reg[31][23]  ( .D(n148), .CP(clk), .Q(\memory[31][23] ) );
  CFD1QXL \memory_reg[31][22]  ( .D(n149), .CP(clk), .Q(\memory[31][22] ) );
  CFD1QXL \memory_reg[31][21]  ( .D(n150), .CP(clk), .Q(\memory[31][21] ) );
  CFD1QXL \memory_reg[31][20]  ( .D(n151), .CP(clk), .Q(\memory[31][20] ) );
  CFD1QXL \memory_reg[31][19]  ( .D(n152), .CP(clk), .Q(\memory[31][19] ) );
  CFD1QXL \memory_reg[31][18]  ( .D(n153), .CP(clk), .Q(\memory[31][18] ) );
  CFD1QXL \memory_reg[31][17]  ( .D(n154), .CP(clk), .Q(\memory[31][17] ) );
  CFD1QXL \memory_reg[31][16]  ( .D(n155), .CP(clk), .Q(\memory[31][16] ) );
  CFD1QXL \memory_reg[31][15]  ( .D(n156), .CP(clk), .Q(\memory[31][15] ) );
  CFD1QXL \memory_reg[31][14]  ( .D(n157), .CP(clk), .Q(\memory[31][14] ) );
  CFD1QXL \memory_reg[31][13]  ( .D(n158), .CP(clk), .Q(\memory[31][13] ) );
  CFD1QXL \memory_reg[31][12]  ( .D(n159), .CP(clk), .Q(\memory[31][12] ) );
  CFD1QXL \memory_reg[31][11]  ( .D(n160), .CP(clk), .Q(\memory[31][11] ) );
  CFD1QXL \memory_reg[31][10]  ( .D(n161), .CP(clk), .Q(\memory[31][10] ) );
  CFD1QXL \memory_reg[31][9]  ( .D(n162), .CP(clk), .Q(\memory[31][9] ) );
  CFD1QXL \memory_reg[31][8]  ( .D(n163), .CP(clk), .Q(\memory[31][8] ) );
  CFD1QXL \memory_reg[31][7]  ( .D(n164), .CP(clk), .Q(\memory[31][7] ) );
  CFD1QXL \memory_reg[31][6]  ( .D(n165), .CP(clk), .Q(\memory[31][6] ) );
  CFD1QXL \memory_reg[31][5]  ( .D(n166), .CP(clk), .Q(\memory[31][5] ) );
  CFD1QXL \memory_reg[31][4]  ( .D(n167), .CP(clk), .Q(\memory[31][4] ) );
  CFD1QXL \memory_reg[31][3]  ( .D(n168), .CP(clk), .Q(\memory[31][3] ) );
  CFD1QXL \memory_reg[31][2]  ( .D(n169), .CP(clk), .Q(\memory[31][2] ) );
  CFD1QXL \memory_reg[31][1]  ( .D(n170), .CP(clk), .Q(\memory[31][1] ) );
  CFD1QXL \memory_reg[31][0]  ( .D(n171), .CP(clk), .Q(\memory[31][0] ) );
  CFD1QXL \memory_reg[7][63]  ( .D(n1812), .CP(clk), .Q(\memory[7][63] ) );
  CFD1QXL \memory_reg[7][62]  ( .D(n1813), .CP(clk), .Q(\memory[7][62] ) );
  CFD1QXL \memory_reg[7][61]  ( .D(n1814), .CP(clk), .Q(\memory[7][61] ) );
  CFD1QXL \memory_reg[7][60]  ( .D(n1815), .CP(clk), .Q(\memory[7][60] ) );
  CFD1QXL \memory_reg[7][59]  ( .D(n1816), .CP(clk), .Q(\memory[7][59] ) );
  CFD1QXL \memory_reg[7][58]  ( .D(n1817), .CP(clk), .Q(\memory[7][58] ) );
  CFD1QXL \memory_reg[7][57]  ( .D(n1818), .CP(clk), .Q(\memory[7][57] ) );
  CFD1QXL \memory_reg[7][56]  ( .D(n1819), .CP(clk), .Q(\memory[7][56] ) );
  CFD1QXL \memory_reg[7][55]  ( .D(n1820), .CP(clk), .Q(\memory[7][55] ) );
  CFD1QXL \memory_reg[7][54]  ( .D(n1821), .CP(clk), .Q(\memory[7][54] ) );
  CFD1QXL \memory_reg[7][53]  ( .D(n1822), .CP(clk), .Q(\memory[7][53] ) );
  CFD1QXL \memory_reg[7][52]  ( .D(n1823), .CP(clk), .Q(\memory[7][52] ) );
  CFD1QXL \memory_reg[7][51]  ( .D(n1824), .CP(clk), .Q(\memory[7][51] ) );
  CFD1QXL \memory_reg[7][50]  ( .D(n1825), .CP(clk), .Q(\memory[7][50] ) );
  CFD1QXL \memory_reg[7][49]  ( .D(n1826), .CP(clk), .Q(\memory[7][49] ) );
  CFD1QXL \memory_reg[7][48]  ( .D(n1827), .CP(clk), .Q(\memory[7][48] ) );
  CFD1QXL \memory_reg[7][47]  ( .D(n1828), .CP(clk), .Q(\memory[7][47] ) );
  CFD1QXL \memory_reg[7][46]  ( .D(n1829), .CP(clk), .Q(\memory[7][46] ) );
  CFD1QXL \memory_reg[7][45]  ( .D(n1830), .CP(clk), .Q(\memory[7][45] ) );
  CFD1QXL \memory_reg[7][44]  ( .D(n1831), .CP(clk), .Q(\memory[7][44] ) );
  CFD1QXL \memory_reg[7][43]  ( .D(n1832), .CP(clk), .Q(\memory[7][43] ) );
  CFD1QXL \memory_reg[7][42]  ( .D(n1833), .CP(clk), .Q(\memory[7][42] ) );
  CFD1QXL \memory_reg[7][41]  ( .D(n1834), .CP(clk), .Q(\memory[7][41] ) );
  CFD1QXL \memory_reg[7][40]  ( .D(n1835), .CP(clk), .Q(\memory[7][40] ) );
  CFD1QXL \memory_reg[7][39]  ( .D(n1836), .CP(clk), .Q(\memory[7][39] ) );
  CFD1QXL \memory_reg[7][38]  ( .D(n1837), .CP(clk), .Q(\memory[7][38] ) );
  CFD1QXL \memory_reg[7][37]  ( .D(n1838), .CP(clk), .Q(\memory[7][37] ) );
  CFD1QXL \memory_reg[7][36]  ( .D(n1839), .CP(clk), .Q(\memory[7][36] ) );
  CFD1QXL \memory_reg[7][35]  ( .D(n1840), .CP(clk), .Q(\memory[7][35] ) );
  CFD1QXL \memory_reg[7][34]  ( .D(n1841), .CP(clk), .Q(\memory[7][34] ) );
  CFD1QXL \memory_reg[7][33]  ( .D(n1842), .CP(clk), .Q(\memory[7][33] ) );
  CFD1QXL \memory_reg[7][32]  ( .D(n1843), .CP(clk), .Q(\memory[7][32] ) );
  CFD1QXL \memory_reg[7][31]  ( .D(n1844), .CP(clk), .Q(\memory[7][31] ) );
  CFD1QXL \memory_reg[7][30]  ( .D(n1845), .CP(clk), .Q(\memory[7][30] ) );
  CFD1QXL \memory_reg[7][29]  ( .D(n1846), .CP(clk), .Q(\memory[7][29] ) );
  CFD1QXL \memory_reg[7][28]  ( .D(n1847), .CP(clk), .Q(\memory[7][28] ) );
  CFD1QXL \memory_reg[7][27]  ( .D(n1848), .CP(clk), .Q(\memory[7][27] ) );
  CFD1QXL \memory_reg[7][26]  ( .D(n1849), .CP(clk), .Q(\memory[7][26] ) );
  CFD1QXL \memory_reg[7][25]  ( .D(n1850), .CP(clk), .Q(\memory[7][25] ) );
  CFD1QXL \memory_reg[7][24]  ( .D(n1851), .CP(clk), .Q(\memory[7][24] ) );
  CFD1QXL \memory_reg[7][23]  ( .D(n1852), .CP(clk), .Q(\memory[7][23] ) );
  CFD1QXL \memory_reg[7][22]  ( .D(n1853), .CP(clk), .Q(\memory[7][22] ) );
  CFD1QXL \memory_reg[7][21]  ( .D(n1854), .CP(clk), .Q(\memory[7][21] ) );
  CFD1QXL \memory_reg[7][20]  ( .D(n1855), .CP(clk), .Q(\memory[7][20] ) );
  CFD1QXL \memory_reg[7][19]  ( .D(n1856), .CP(clk), .Q(\memory[7][19] ) );
  CFD1QXL \memory_reg[7][18]  ( .D(n1857), .CP(clk), .Q(\memory[7][18] ) );
  CFD1QXL \memory_reg[7][17]  ( .D(n1858), .CP(clk), .Q(\memory[7][17] ) );
  CFD1QXL \memory_reg[7][16]  ( .D(n1859), .CP(clk), .Q(\memory[7][16] ) );
  CFD1QXL \memory_reg[7][15]  ( .D(n1860), .CP(clk), .Q(\memory[7][15] ) );
  CFD1QXL \memory_reg[7][14]  ( .D(n1861), .CP(clk), .Q(\memory[7][14] ) );
  CFD1QXL \memory_reg[7][13]  ( .D(n1862), .CP(clk), .Q(\memory[7][13] ) );
  CFD1QXL \memory_reg[7][12]  ( .D(n1863), .CP(clk), .Q(\memory[7][12] ) );
  CFD1QXL \memory_reg[7][11]  ( .D(n1864), .CP(clk), .Q(\memory[7][11] ) );
  CFD1QXL \memory_reg[7][10]  ( .D(n1865), .CP(clk), .Q(\memory[7][10] ) );
  CFD1QXL \memory_reg[7][9]  ( .D(n1866), .CP(clk), .Q(\memory[7][9] ) );
  CFD1QXL \memory_reg[7][8]  ( .D(n1867), .CP(clk), .Q(\memory[7][8] ) );
  CFD1QXL \memory_reg[7][7]  ( .D(n1868), .CP(clk), .Q(\memory[7][7] ) );
  CFD1QXL \memory_reg[7][6]  ( .D(n1869), .CP(clk), .Q(\memory[7][6] ) );
  CFD1QXL \memory_reg[7][5]  ( .D(n1870), .CP(clk), .Q(\memory[7][5] ) );
  CFD1QXL \memory_reg[7][4]  ( .D(n1871), .CP(clk), .Q(\memory[7][4] ) );
  CFD1QXL \memory_reg[7][3]  ( .D(n1872), .CP(clk), .Q(\memory[7][3] ) );
  CFD1QXL \memory_reg[7][2]  ( .D(n1873), .CP(clk), .Q(\memory[7][2] ) );
  CFD1QXL \memory_reg[7][1]  ( .D(n1874), .CP(clk), .Q(\memory[7][1] ) );
  CFD1QXL \memory_reg[7][0]  ( .D(n1875), .CP(clk), .Q(\memory[7][0] ) );
  CFD1QXL \lenout_reg[5]  ( .D(n2452), .CP(clk), .Q(lenout[5]) );
  CFD1QXL \lenout_reg[6]  ( .D(n2453), .CP(clk), .Q(lenout[6]) );
  CFD1QXL \lenout_reg[4]  ( .D(n2451), .CP(clk), .Q(lenout[4]) );
  CFD1QXL \lenout_reg[3]  ( .D(n2450), .CP(clk), .Q(lenout[3]) );
  CFD1QXL \lenout_reg[2]  ( .D(n2449), .CP(clk), .Q(lenout[2]) );
  CFD1QXL \lenout_reg[1]  ( .D(n2448), .CP(clk), .Q(lenout[1]) );
  CFD1QXL \lenout_reg[0]  ( .D(n2447), .CP(clk), .Q(lenout[0]) );
  CFD1QXL \dataout_reg[63]  ( .D(n2446), .CP(clk), .Q(dataout[63]) );
  CFD1QXL \dataout_reg[62]  ( .D(n2445), .CP(clk), .Q(dataout[62]) );
  CFD1QXL \dataout_reg[61]  ( .D(n2444), .CP(clk), .Q(dataout[61]) );
  CFD1QXL \dataout_reg[60]  ( .D(n2443), .CP(clk), .Q(dataout[60]) );
  CFD1QXL \dataout_reg[59]  ( .D(n2442), .CP(clk), .Q(dataout[59]) );
  CFD1QXL \dataout_reg[58]  ( .D(n2441), .CP(clk), .Q(dataout[58]) );
  CFD1QXL \dataout_reg[57]  ( .D(n2440), .CP(clk), .Q(dataout[57]) );
  CFD1QXL \dataout_reg[56]  ( .D(n2439), .CP(clk), .Q(dataout[56]) );
  CFD1QXL \dataout_reg[55]  ( .D(n2438), .CP(clk), .Q(dataout[55]) );
  CFD1QXL \dataout_reg[54]  ( .D(n2437), .CP(clk), .Q(dataout[54]) );
  CFD1QXL \dataout_reg[53]  ( .D(n2436), .CP(clk), .Q(dataout[53]) );
  CFD1QXL \dataout_reg[52]  ( .D(n2435), .CP(clk), .Q(dataout[52]) );
  CFD1QXL \dataout_reg[51]  ( .D(n2434), .CP(clk), .Q(dataout[51]) );
  CFD1QXL \dataout_reg[50]  ( .D(n2433), .CP(clk), .Q(dataout[50]) );
  CFD1QXL \dataout_reg[49]  ( .D(n2432), .CP(clk), .Q(dataout[49]) );
  CFD1QXL \dataout_reg[48]  ( .D(n2431), .CP(clk), .Q(dataout[48]) );
  CFD1QXL \dataout_reg[47]  ( .D(n2430), .CP(clk), .Q(dataout[47]) );
  CFD1QXL \dataout_reg[46]  ( .D(n2429), .CP(clk), .Q(dataout[46]) );
  CFD1QXL \dataout_reg[45]  ( .D(n2428), .CP(clk), .Q(dataout[45]) );
  CFD1QXL \dataout_reg[44]  ( .D(n2427), .CP(clk), .Q(dataout[44]) );
  CFD1QXL \dataout_reg[43]  ( .D(n2426), .CP(clk), .Q(dataout[43]) );
  CFD1QXL \dataout_reg[42]  ( .D(n2425), .CP(clk), .Q(dataout[42]) );
  CFD1QXL \dataout_reg[41]  ( .D(n2424), .CP(clk), .Q(dataout[41]) );
  CFD1QXL \dataout_reg[40]  ( .D(n2423), .CP(clk), .Q(dataout[40]) );
  CFD1QXL \dataout_reg[39]  ( .D(n2422), .CP(clk), .Q(dataout[39]) );
  CFD1QXL \dataout_reg[38]  ( .D(n2421), .CP(clk), .Q(dataout[38]) );
  CFD1QXL \dataout_reg[37]  ( .D(n2420), .CP(clk), .Q(dataout[37]) );
  CFD1QXL \dataout_reg[36]  ( .D(n2419), .CP(clk), .Q(dataout[36]) );
  CFD1QXL \dataout_reg[35]  ( .D(n2418), .CP(clk), .Q(dataout[35]) );
  CFD1QXL \dataout_reg[34]  ( .D(n2417), .CP(clk), .Q(dataout[34]) );
  CFD1QXL \dataout_reg[33]  ( .D(n2416), .CP(clk), .Q(dataout[33]) );
  CFD1QXL \dataout_reg[32]  ( .D(n2415), .CP(clk), .Q(dataout[32]) );
  CFD1QXL \dataout_reg[31]  ( .D(n2414), .CP(clk), .Q(dataout[31]) );
  CFD1QXL \dataout_reg[30]  ( .D(n2413), .CP(clk), .Q(dataout[30]) );
  CFD1QXL \dataout_reg[29]  ( .D(n2412), .CP(clk), .Q(dataout[29]) );
  CFD1QXL \dataout_reg[28]  ( .D(n2411), .CP(clk), .Q(dataout[28]) );
  CFD1QXL \dataout_reg[27]  ( .D(n2410), .CP(clk), .Q(dataout[27]) );
  CFD1QXL \dataout_reg[26]  ( .D(n2409), .CP(clk), .Q(dataout[26]) );
  CFD1QXL \dataout_reg[25]  ( .D(n2408), .CP(clk), .Q(dataout[25]) );
  CFD1QXL \dataout_reg[24]  ( .D(n2407), .CP(clk), .Q(dataout[24]) );
  CFD1QXL \dataout_reg[23]  ( .D(n2406), .CP(clk), .Q(dataout[23]) );
  CFD1QXL \dataout_reg[22]  ( .D(n2405), .CP(clk), .Q(dataout[22]) );
  CFD1QXL \dataout_reg[21]  ( .D(n2404), .CP(clk), .Q(dataout[21]) );
  CFD1QXL \dataout_reg[20]  ( .D(n2403), .CP(clk), .Q(dataout[20]) );
  CFD1QXL \dataout_reg[19]  ( .D(n2402), .CP(clk), .Q(dataout[19]) );
  CFD1QXL \dataout_reg[18]  ( .D(n2401), .CP(clk), .Q(dataout[18]) );
  CFD1QXL \dataout_reg[17]  ( .D(n2400), .CP(clk), .Q(dataout[17]) );
  CFD1QXL \dataout_reg[16]  ( .D(n2399), .CP(clk), .Q(dataout[16]) );
  CFD1QXL \dataout_reg[15]  ( .D(n2398), .CP(clk), .Q(dataout[15]) );
  CFD1QXL \dataout_reg[14]  ( .D(n2397), .CP(clk), .Q(dataout[14]) );
  CFD1QXL \dataout_reg[13]  ( .D(n2396), .CP(clk), .Q(dataout[13]) );
  CFD1QXL \dataout_reg[12]  ( .D(n2395), .CP(clk), .Q(dataout[12]) );
  CFD1QXL \dataout_reg[11]  ( .D(n2394), .CP(clk), .Q(dataout[11]) );
  CFD1QXL \dataout_reg[10]  ( .D(n2393), .CP(clk), .Q(dataout[10]) );
  CFD1QXL \dataout_reg[9]  ( .D(n2392), .CP(clk), .Q(dataout[9]) );
  CFD1QXL \dataout_reg[8]  ( .D(n2391), .CP(clk), .Q(dataout[8]) );
  CFD1QXL \dataout_reg[7]  ( .D(n2390), .CP(clk), .Q(dataout[7]) );
  CFD1QXL \dataout_reg[6]  ( .D(n2389), .CP(clk), .Q(dataout[6]) );
  CFD1QXL \dataout_reg[5]  ( .D(n2388), .CP(clk), .Q(dataout[5]) );
  CFD1QXL \dataout_reg[4]  ( .D(n2387), .CP(clk), .Q(dataout[4]) );
  CFD1QXL \dataout_reg[3]  ( .D(n2386), .CP(clk), .Q(dataout[3]) );
  CFD1QXL \dataout_reg[2]  ( .D(n2385), .CP(clk), .Q(dataout[2]) );
  CFD1QXL \dataout_reg[1]  ( .D(n2384), .CP(clk), .Q(dataout[1]) );
  CFD1QXL \dataout_reg[0]  ( .D(n2383), .CP(clk), .Q(dataout[0]) );
  CFD1QXL \memory_reg[27][62]  ( .D(n393), .CP(clk), .Q(\memory[27][62] ) );
  CFD1QXL \memory_reg[23][62]  ( .D(n677), .CP(clk), .Q(\memory[23][62] ) );
  CFD1QXL \memory_reg[19][62]  ( .D(n961), .CP(clk), .Q(\memory[19][62] ) );
  CFD1QXL \memory_reg[15][62]  ( .D(n1245), .CP(clk), .Q(\memory[15][62] ) );
  CFD1QXL \out_new_reg[63]  ( .D(n76), .CP(clk), .Q(out_new[63]) );
  CFD1QXL \out_new_reg[62]  ( .D(n75), .CP(clk), .Q(out_new[62]) );
  CFD1QXL \out_new_reg[61]  ( .D(n74), .CP(clk), .Q(out_new[61]) );
  CFD1QXL \out_new_reg[60]  ( .D(n73), .CP(clk), .Q(out_new[60]) );
  CFD1QXL \out_new_reg[59]  ( .D(n72), .CP(clk), .Q(out_new[59]) );
  CFD1QXL \out_new_reg[58]  ( .D(n71), .CP(clk), .Q(out_new[58]) );
  CFD1QXL \out_new_reg[57]  ( .D(n70), .CP(clk), .Q(out_new[57]) );
  CFD1QXL \out_new_reg[56]  ( .D(n69), .CP(clk), .Q(out_new[56]) );
  CFD1QXL \out_new_reg[55]  ( .D(n68), .CP(clk), .Q(out_new[55]) );
  CFD1QXL \out_new_reg[54]  ( .D(n67), .CP(clk), .Q(out_new[54]) );
  CFD1QXL \out_new_reg[53]  ( .D(n66), .CP(clk), .Q(out_new[53]) );
  CFD1QXL \out_new_reg[52]  ( .D(n65), .CP(clk), .Q(out_new[52]) );
  CFD1QXL \out_new_reg[51]  ( .D(n64), .CP(clk), .Q(out_new[51]) );
  CFD1QXL \out_new_reg[50]  ( .D(n63), .CP(clk), .Q(out_new[50]) );
  CFD1QXL \out_new_reg[49]  ( .D(n62), .CP(clk), .Q(out_new[49]) );
  CFD1QXL \out_new_reg[48]  ( .D(n61), .CP(clk), .Q(out_new[48]) );
  CFD1QXL \out_new_reg[47]  ( .D(n60), .CP(clk), .Q(out_new[47]) );
  CFD1QXL \out_new_reg[46]  ( .D(n59), .CP(clk), .Q(out_new[46]) );
  CFD1QXL \out_new_reg[45]  ( .D(n58), .CP(clk), .Q(out_new[45]) );
  CFD1QXL \out_new_reg[44]  ( .D(n57), .CP(clk), .Q(out_new[44]) );
  CFD1QXL \out_new_reg[43]  ( .D(n56), .CP(clk), .Q(out_new[43]) );
  CFD1QXL \out_new_reg[42]  ( .D(n55), .CP(clk), .Q(out_new[42]) );
  CFD1QXL \out_new_reg[41]  ( .D(n54), .CP(clk), .Q(out_new[41]) );
  CFD1QXL \out_new_reg[40]  ( .D(n53), .CP(clk), .Q(out_new[40]) );
  CFD1QXL \out_new_reg[39]  ( .D(n52), .CP(clk), .Q(out_new[39]) );
  CFD1QXL \out_new_reg[38]  ( .D(n51), .CP(clk), .Q(out_new[38]) );
  CFD1QXL \out_new_reg[37]  ( .D(n50), .CP(clk), .Q(out_new[37]) );
  CFD1QXL \out_new_reg[36]  ( .D(n49), .CP(clk), .Q(out_new[36]) );
  CFD1QXL \out_new_reg[35]  ( .D(n48), .CP(clk), .Q(out_new[35]) );
  CFD1QXL \out_new_reg[34]  ( .D(n47), .CP(clk), .Q(out_new[34]) );
  CFD1QXL \out_new_reg[33]  ( .D(n46), .CP(clk), .Q(out_new[33]) );
  CFD1QXL \out_new_reg[32]  ( .D(n45), .CP(clk), .Q(out_new[32]) );
  CFD1QXL \out_new_reg[31]  ( .D(n44), .CP(clk), .Q(out_new[31]) );
  CFD1QXL \out_new_reg[30]  ( .D(n43), .CP(clk), .Q(out_new[30]) );
  CFD1QXL \out_new_reg[29]  ( .D(n42), .CP(clk), .Q(out_new[29]) );
  CFD1QXL \out_new_reg[28]  ( .D(n41), .CP(clk), .Q(out_new[28]) );
  CFD1QXL \out_new_reg[27]  ( .D(n40), .CP(clk), .Q(out_new[27]) );
  CFD1QXL \out_new_reg[26]  ( .D(n39), .CP(clk), .Q(out_new[26]) );
  CFD1QXL \out_new_reg[25]  ( .D(n38), .CP(clk), .Q(out_new[25]) );
  CFD1QXL \out_new_reg[24]  ( .D(n37), .CP(clk), .Q(out_new[24]) );
  CFD1QXL \out_new_reg[23]  ( .D(n36), .CP(clk), .Q(out_new[23]) );
  CFD1QXL \out_new_reg[22]  ( .D(n35), .CP(clk), .Q(out_new[22]) );
  CFD1QXL \out_new_reg[21]  ( .D(n34), .CP(clk), .Q(out_new[21]) );
  CFD1QXL \out_new_reg[20]  ( .D(n33), .CP(clk), .Q(out_new[20]) );
  CFD1QXL \out_new_reg[19]  ( .D(n32), .CP(clk), .Q(out_new[19]) );
  CFD1QXL \out_new_reg[18]  ( .D(n31), .CP(clk), .Q(out_new[18]) );
  CFD1QXL \out_new_reg[17]  ( .D(n30), .CP(clk), .Q(out_new[17]) );
  CFD1QXL \out_new_reg[16]  ( .D(n29), .CP(clk), .Q(out_new[16]) );
  CFD1QXL \out_new_reg[15]  ( .D(n28), .CP(clk), .Q(out_new[15]) );
  CFD1QXL \out_new_reg[14]  ( .D(n27), .CP(clk), .Q(out_new[14]) );
  CFD1QXL \out_new_reg[13]  ( .D(n26), .CP(clk), .Q(out_new[13]) );
  CFD1QXL \out_new_reg[12]  ( .D(n25), .CP(clk), .Q(out_new[12]) );
  CFD1QXL \out_new_reg[11]  ( .D(n24), .CP(clk), .Q(out_new[11]) );
  CFD1QXL \out_new_reg[10]  ( .D(n23), .CP(clk), .Q(out_new[10]) );
  CFD1QXL \out_new_reg[9]  ( .D(n22), .CP(clk), .Q(out_new[9]) );
  CFD1QXL \out_new_reg[8]  ( .D(n21), .CP(clk), .Q(out_new[8]) );
  CFD1QXL \out_new_reg[7]  ( .D(n20), .CP(clk), .Q(out_new[7]) );
  CFD1QXL \out_new_reg[6]  ( .D(n19), .CP(clk), .Q(out_new[6]) );
  CFD1QXL \out_new_reg[5]  ( .D(n18), .CP(clk), .Q(out_new[5]) );
  CFD1QXL \out_new_reg[4]  ( .D(n17), .CP(clk), .Q(out_new[4]) );
  CFD1QXL \out_new_reg[3]  ( .D(n16), .CP(clk), .Q(out_new[3]) );
  CFD1QXL \out_new_reg[2]  ( .D(n15), .CP(clk), .Q(out_new[2]) );
  CFD1QXL \out_new_reg[1]  ( .D(n14), .CP(clk), .Q(out_new[1]) );
  CFD1QXL \out_new_reg[0]  ( .D(n13), .CP(clk), .Q(out_new[0]) );
  CFD1QXL \lout_new_reg[6]  ( .D(n6), .CP(clk), .Q(lout_new[6]) );
  CFD1QXL \lout_new_reg[5]  ( .D(n7), .CP(clk), .Q(lout_new[5]) );
  CFD1QXL \lout_new_reg[4]  ( .D(n8), .CP(clk), .Q(lout_new[4]) );
  CFD1QXL \lout_new_reg[3]  ( .D(n9), .CP(clk), .Q(lout_new[3]) );
  CFD1QXL \lout_new_reg[2]  ( .D(n10), .CP(clk), .Q(lout_new[2]) );
  CFD1QXL \lout_new_reg[1]  ( .D(n11), .CP(clk), .Q(lout_new[1]) );
  CFD1QXL \lout_new_reg[0]  ( .D(n12), .CP(clk), .Q(lout_new[0]) );
  CFD1QXL \memory_reg[27][63]  ( .D(n392), .CP(clk), .Q(\memory[27][63] ) );
  CFD1QXL \memory_reg[27][61]  ( .D(n394), .CP(clk), .Q(\memory[27][61] ) );
  CFD1QXL \memory_reg[27][60]  ( .D(n395), .CP(clk), .Q(\memory[27][60] ) );
  CFD1QXL \memory_reg[27][59]  ( .D(n396), .CP(clk), .Q(\memory[27][59] ) );
  CFD1QXL \memory_reg[27][58]  ( .D(n397), .CP(clk), .Q(\memory[27][58] ) );
  CFD1QXL \memory_reg[27][57]  ( .D(n398), .CP(clk), .Q(\memory[27][57] ) );
  CFD1QXL \memory_reg[27][56]  ( .D(n399), .CP(clk), .Q(\memory[27][56] ) );
  CFD1QXL \memory_reg[27][55]  ( .D(n400), .CP(clk), .Q(\memory[27][55] ) );
  CFD1QXL \memory_reg[27][54]  ( .D(n401), .CP(clk), .Q(\memory[27][54] ) );
  CFD1QXL \memory_reg[27][53]  ( .D(n402), .CP(clk), .Q(\memory[27][53] ) );
  CFD1QXL \memory_reg[27][52]  ( .D(n403), .CP(clk), .Q(\memory[27][52] ) );
  CFD1QXL \memory_reg[27][51]  ( .D(n404), .CP(clk), .Q(\memory[27][51] ) );
  CFD1QXL \memory_reg[27][50]  ( .D(n405), .CP(clk), .Q(\memory[27][50] ) );
  CFD1QXL \memory_reg[27][49]  ( .D(n406), .CP(clk), .Q(\memory[27][49] ) );
  CFD1QXL \memory_reg[27][48]  ( .D(n407), .CP(clk), .Q(\memory[27][48] ) );
  CFD1QXL \memory_reg[27][47]  ( .D(n408), .CP(clk), .Q(\memory[27][47] ) );
  CFD1QXL \memory_reg[27][46]  ( .D(n409), .CP(clk), .Q(\memory[27][46] ) );
  CFD1QXL \memory_reg[27][45]  ( .D(n410), .CP(clk), .Q(\memory[27][45] ) );
  CFD1QXL \memory_reg[27][44]  ( .D(n411), .CP(clk), .Q(\memory[27][44] ) );
  CFD1QXL \memory_reg[27][43]  ( .D(n412), .CP(clk), .Q(\memory[27][43] ) );
  CFD1QXL \memory_reg[27][42]  ( .D(n413), .CP(clk), .Q(\memory[27][42] ) );
  CFD1QXL \memory_reg[27][41]  ( .D(n414), .CP(clk), .Q(\memory[27][41] ) );
  CFD1QXL \memory_reg[27][40]  ( .D(n415), .CP(clk), .Q(\memory[27][40] ) );
  CFD1QXL \memory_reg[27][39]  ( .D(n416), .CP(clk), .Q(\memory[27][39] ) );
  CFD1QXL \memory_reg[27][38]  ( .D(n417), .CP(clk), .Q(\memory[27][38] ) );
  CFD1QXL \memory_reg[27][37]  ( .D(n418), .CP(clk), .Q(\memory[27][37] ) );
  CFD1QXL \memory_reg[27][36]  ( .D(n419), .CP(clk), .Q(\memory[27][36] ) );
  CFD1QXL \memory_reg[27][35]  ( .D(n420), .CP(clk), .Q(\memory[27][35] ) );
  CFD1QXL \memory_reg[27][34]  ( .D(n421), .CP(clk), .Q(\memory[27][34] ) );
  CFD1QXL \memory_reg[27][33]  ( .D(n422), .CP(clk), .Q(\memory[27][33] ) );
  CFD1QXL \memory_reg[27][32]  ( .D(n423), .CP(clk), .Q(\memory[27][32] ) );
  CFD1QXL \memory_reg[27][31]  ( .D(n424), .CP(clk), .Q(\memory[27][31] ) );
  CFD1QXL \memory_reg[27][30]  ( .D(n425), .CP(clk), .Q(\memory[27][30] ) );
  CFD1QXL \memory_reg[27][29]  ( .D(n426), .CP(clk), .Q(\memory[27][29] ) );
  CFD1QXL \memory_reg[27][28]  ( .D(n427), .CP(clk), .Q(\memory[27][28] ) );
  CFD1QXL \memory_reg[27][27]  ( .D(n428), .CP(clk), .Q(\memory[27][27] ) );
  CFD1QXL \memory_reg[27][26]  ( .D(n429), .CP(clk), .Q(\memory[27][26] ) );
  CFD1QXL \memory_reg[27][25]  ( .D(n430), .CP(clk), .Q(\memory[27][25] ) );
  CFD1QXL \memory_reg[27][24]  ( .D(n431), .CP(clk), .Q(\memory[27][24] ) );
  CFD1QXL \memory_reg[27][23]  ( .D(n432), .CP(clk), .Q(\memory[27][23] ) );
  CFD1QXL \memory_reg[27][22]  ( .D(n433), .CP(clk), .Q(\memory[27][22] ) );
  CFD1QXL \memory_reg[27][21]  ( .D(n434), .CP(clk), .Q(\memory[27][21] ) );
  CFD1QXL \memory_reg[27][20]  ( .D(n435), .CP(clk), .Q(\memory[27][20] ) );
  CFD1QXL \memory_reg[27][19]  ( .D(n436), .CP(clk), .Q(\memory[27][19] ) );
  CFD1QXL \memory_reg[27][18]  ( .D(n437), .CP(clk), .Q(\memory[27][18] ) );
  CFD1QXL \memory_reg[27][17]  ( .D(n438), .CP(clk), .Q(\memory[27][17] ) );
  CFD1QXL \memory_reg[27][16]  ( .D(n439), .CP(clk), .Q(\memory[27][16] ) );
  CFD1QXL \memory_reg[27][15]  ( .D(n440), .CP(clk), .Q(\memory[27][15] ) );
  CFD1QXL \memory_reg[27][14]  ( .D(n441), .CP(clk), .Q(\memory[27][14] ) );
  CFD1QXL \memory_reg[27][13]  ( .D(n442), .CP(clk), .Q(\memory[27][13] ) );
  CFD1QXL \memory_reg[27][12]  ( .D(n443), .CP(clk), .Q(\memory[27][12] ) );
  CFD1QXL \memory_reg[27][11]  ( .D(n444), .CP(clk), .Q(\memory[27][11] ) );
  CFD1QXL \memory_reg[27][10]  ( .D(n445), .CP(clk), .Q(\memory[27][10] ) );
  CFD1QXL \memory_reg[27][9]  ( .D(n446), .CP(clk), .Q(\memory[27][9] ) );
  CFD1QXL \memory_reg[27][8]  ( .D(n447), .CP(clk), .Q(\memory[27][8] ) );
  CFD1QXL \memory_reg[27][7]  ( .D(n448), .CP(clk), .Q(\memory[27][7] ) );
  CFD1QXL \memory_reg[27][6]  ( .D(n449), .CP(clk), .Q(\memory[27][6] ) );
  CFD1QXL \memory_reg[27][5]  ( .D(n450), .CP(clk), .Q(\memory[27][5] ) );
  CFD1QXL \memory_reg[27][4]  ( .D(n451), .CP(clk), .Q(\memory[27][4] ) );
  CFD1QXL \memory_reg[27][3]  ( .D(n452), .CP(clk), .Q(\memory[27][3] ) );
  CFD1QXL \memory_reg[27][2]  ( .D(n453), .CP(clk), .Q(\memory[27][2] ) );
  CFD1QXL \memory_reg[27][1]  ( .D(n454), .CP(clk), .Q(\memory[27][1] ) );
  CFD1QXL \memory_reg[27][0]  ( .D(n455), .CP(clk), .Q(\memory[27][0] ) );
  CFD1QXL \memory_reg[23][63]  ( .D(n676), .CP(clk), .Q(\memory[23][63] ) );
  CFD1QXL \memory_reg[23][61]  ( .D(n678), .CP(clk), .Q(\memory[23][61] ) );
  CFD1QXL \memory_reg[23][60]  ( .D(n679), .CP(clk), .Q(\memory[23][60] ) );
  CFD1QXL \memory_reg[23][59]  ( .D(n680), .CP(clk), .Q(\memory[23][59] ) );
  CFD1QXL \memory_reg[23][58]  ( .D(n681), .CP(clk), .Q(\memory[23][58] ) );
  CFD1QXL \memory_reg[23][57]  ( .D(n682), .CP(clk), .Q(\memory[23][57] ) );
  CFD1QXL \memory_reg[23][56]  ( .D(n683), .CP(clk), .Q(\memory[23][56] ) );
  CFD1QXL \memory_reg[23][55]  ( .D(n684), .CP(clk), .Q(\memory[23][55] ) );
  CFD1QXL \memory_reg[23][54]  ( .D(n685), .CP(clk), .Q(\memory[23][54] ) );
  CFD1QXL \memory_reg[23][53]  ( .D(n686), .CP(clk), .Q(\memory[23][53] ) );
  CFD1QXL \memory_reg[23][52]  ( .D(n687), .CP(clk), .Q(\memory[23][52] ) );
  CFD1QXL \memory_reg[23][51]  ( .D(n688), .CP(clk), .Q(\memory[23][51] ) );
  CFD1QXL \memory_reg[23][50]  ( .D(n689), .CP(clk), .Q(\memory[23][50] ) );
  CFD1QXL \memory_reg[23][49]  ( .D(n690), .CP(clk), .Q(\memory[23][49] ) );
  CFD1QXL \memory_reg[23][48]  ( .D(n691), .CP(clk), .Q(\memory[23][48] ) );
  CFD1QXL \memory_reg[23][47]  ( .D(n692), .CP(clk), .Q(\memory[23][47] ) );
  CFD1QXL \memory_reg[23][46]  ( .D(n693), .CP(clk), .Q(\memory[23][46] ) );
  CFD1QXL \memory_reg[23][45]  ( .D(n694), .CP(clk), .Q(\memory[23][45] ) );
  CFD1QXL \memory_reg[23][44]  ( .D(n695), .CP(clk), .Q(\memory[23][44] ) );
  CFD1QXL \memory_reg[23][43]  ( .D(n696), .CP(clk), .Q(\memory[23][43] ) );
  CFD1QXL \memory_reg[23][42]  ( .D(n697), .CP(clk), .Q(\memory[23][42] ) );
  CFD1QXL \memory_reg[23][41]  ( .D(n698), .CP(clk), .Q(\memory[23][41] ) );
  CFD1QXL \memory_reg[23][40]  ( .D(n699), .CP(clk), .Q(\memory[23][40] ) );
  CFD1QXL \memory_reg[23][39]  ( .D(n700), .CP(clk), .Q(\memory[23][39] ) );
  CFD1QXL \memory_reg[23][38]  ( .D(n701), .CP(clk), .Q(\memory[23][38] ) );
  CFD1QXL \memory_reg[23][37]  ( .D(n702), .CP(clk), .Q(\memory[23][37] ) );
  CFD1QXL \memory_reg[23][36]  ( .D(n703), .CP(clk), .Q(\memory[23][36] ) );
  CFD1QXL \memory_reg[23][35]  ( .D(n704), .CP(clk), .Q(\memory[23][35] ) );
  CFD1QXL \memory_reg[23][34]  ( .D(n705), .CP(clk), .Q(\memory[23][34] ) );
  CFD1QXL \memory_reg[23][33]  ( .D(n706), .CP(clk), .Q(\memory[23][33] ) );
  CFD1QXL \memory_reg[23][32]  ( .D(n707), .CP(clk), .Q(\memory[23][32] ) );
  CFD1QXL \memory_reg[23][31]  ( .D(n708), .CP(clk), .Q(\memory[23][31] ) );
  CFD1QXL \memory_reg[23][30]  ( .D(n709), .CP(clk), .Q(\memory[23][30] ) );
  CFD1QXL \memory_reg[23][29]  ( .D(n710), .CP(clk), .Q(\memory[23][29] ) );
  CFD1QXL \memory_reg[23][28]  ( .D(n711), .CP(clk), .Q(\memory[23][28] ) );
  CFD1QXL \memory_reg[23][27]  ( .D(n712), .CP(clk), .Q(\memory[23][27] ) );
  CFD1QXL \memory_reg[23][26]  ( .D(n713), .CP(clk), .Q(\memory[23][26] ) );
  CFD1QXL \memory_reg[23][25]  ( .D(n714), .CP(clk), .Q(\memory[23][25] ) );
  CFD1QXL \memory_reg[23][24]  ( .D(n715), .CP(clk), .Q(\memory[23][24] ) );
  CFD1QXL \memory_reg[23][23]  ( .D(n716), .CP(clk), .Q(\memory[23][23] ) );
  CFD1QXL \memory_reg[23][22]  ( .D(n717), .CP(clk), .Q(\memory[23][22] ) );
  CFD1QXL \memory_reg[23][21]  ( .D(n718), .CP(clk), .Q(\memory[23][21] ) );
  CFD1QXL \memory_reg[23][20]  ( .D(n719), .CP(clk), .Q(\memory[23][20] ) );
  CFD1QXL \memory_reg[23][19]  ( .D(n720), .CP(clk), .Q(\memory[23][19] ) );
  CFD1QXL \memory_reg[23][18]  ( .D(n721), .CP(clk), .Q(\memory[23][18] ) );
  CFD1QXL \memory_reg[23][17]  ( .D(n722), .CP(clk), .Q(\memory[23][17] ) );
  CFD1QXL \memory_reg[23][16]  ( .D(n723), .CP(clk), .Q(\memory[23][16] ) );
  CFD1QXL \memory_reg[23][15]  ( .D(n724), .CP(clk), .Q(\memory[23][15] ) );
  CFD1QXL \memory_reg[23][14]  ( .D(n725), .CP(clk), .Q(\memory[23][14] ) );
  CFD1QXL \memory_reg[23][13]  ( .D(n726), .CP(clk), .Q(\memory[23][13] ) );
  CFD1QXL \memory_reg[23][12]  ( .D(n727), .CP(clk), .Q(\memory[23][12] ) );
  CFD1QXL \memory_reg[23][11]  ( .D(n728), .CP(clk), .Q(\memory[23][11] ) );
  CFD1QXL \memory_reg[23][10]  ( .D(n729), .CP(clk), .Q(\memory[23][10] ) );
  CFD1QXL \memory_reg[23][9]  ( .D(n730), .CP(clk), .Q(\memory[23][9] ) );
  CFD1QXL \memory_reg[23][8]  ( .D(n731), .CP(clk), .Q(\memory[23][8] ) );
  CFD1QXL \memory_reg[23][7]  ( .D(n732), .CP(clk), .Q(\memory[23][7] ) );
  CFD1QXL \memory_reg[23][6]  ( .D(n733), .CP(clk), .Q(\memory[23][6] ) );
  CFD1QXL \memory_reg[23][5]  ( .D(n734), .CP(clk), .Q(\memory[23][5] ) );
  CFD1QXL \memory_reg[23][4]  ( .D(n735), .CP(clk), .Q(\memory[23][4] ) );
  CFD1QXL \memory_reg[23][3]  ( .D(n736), .CP(clk), .Q(\memory[23][3] ) );
  CFD1QXL \memory_reg[23][2]  ( .D(n737), .CP(clk), .Q(\memory[23][2] ) );
  CFD1QXL \memory_reg[23][1]  ( .D(n738), .CP(clk), .Q(\memory[23][1] ) );
  CFD1QXL \memory_reg[23][0]  ( .D(n739), .CP(clk), .Q(\memory[23][0] ) );
  CFD1QXL \memory_reg[19][63]  ( .D(n960), .CP(clk), .Q(\memory[19][63] ) );
  CFD1QXL \memory_reg[19][61]  ( .D(n962), .CP(clk), .Q(\memory[19][61] ) );
  CFD1QXL \memory_reg[19][60]  ( .D(n963), .CP(clk), .Q(\memory[19][60] ) );
  CFD1QXL \memory_reg[19][59]  ( .D(n964), .CP(clk), .Q(\memory[19][59] ) );
  CFD1QXL \memory_reg[19][58]  ( .D(n965), .CP(clk), .Q(\memory[19][58] ) );
  CFD1QXL \memory_reg[19][57]  ( .D(n966), .CP(clk), .Q(\memory[19][57] ) );
  CFD1QXL \memory_reg[19][56]  ( .D(n967), .CP(clk), .Q(\memory[19][56] ) );
  CFD1QXL \memory_reg[19][55]  ( .D(n968), .CP(clk), .Q(\memory[19][55] ) );
  CFD1QXL \memory_reg[19][54]  ( .D(n969), .CP(clk), .Q(\memory[19][54] ) );
  CFD1QXL \memory_reg[19][53]  ( .D(n970), .CP(clk), .Q(\memory[19][53] ) );
  CFD1QXL \memory_reg[19][52]  ( .D(n971), .CP(clk), .Q(\memory[19][52] ) );
  CFD1QXL \memory_reg[19][51]  ( .D(n972), .CP(clk), .Q(\memory[19][51] ) );
  CFD1QXL \memory_reg[19][50]  ( .D(n973), .CP(clk), .Q(\memory[19][50] ) );
  CFD1QXL \memory_reg[19][49]  ( .D(n974), .CP(clk), .Q(\memory[19][49] ) );
  CFD1QXL \memory_reg[19][48]  ( .D(n975), .CP(clk), .Q(\memory[19][48] ) );
  CFD1QXL \memory_reg[19][47]  ( .D(n976), .CP(clk), .Q(\memory[19][47] ) );
  CFD1QXL \memory_reg[19][46]  ( .D(n977), .CP(clk), .Q(\memory[19][46] ) );
  CFD1QXL \memory_reg[19][45]  ( .D(n978), .CP(clk), .Q(\memory[19][45] ) );
  CFD1QXL \memory_reg[19][44]  ( .D(n979), .CP(clk), .Q(\memory[19][44] ) );
  CFD1QXL \memory_reg[19][43]  ( .D(n980), .CP(clk), .Q(\memory[19][43] ) );
  CFD1QXL \memory_reg[19][42]  ( .D(n981), .CP(clk), .Q(\memory[19][42] ) );
  CFD1QXL \memory_reg[19][41]  ( .D(n982), .CP(clk), .Q(\memory[19][41] ) );
  CFD1QXL \memory_reg[19][40]  ( .D(n983), .CP(clk), .Q(\memory[19][40] ) );
  CFD1QXL \memory_reg[19][39]  ( .D(n984), .CP(clk), .Q(\memory[19][39] ) );
  CFD1QXL \memory_reg[19][38]  ( .D(n985), .CP(clk), .Q(\memory[19][38] ) );
  CFD1QXL \memory_reg[19][37]  ( .D(n986), .CP(clk), .Q(\memory[19][37] ) );
  CFD1QXL \memory_reg[19][36]  ( .D(n987), .CP(clk), .Q(\memory[19][36] ) );
  CFD1QXL \memory_reg[19][35]  ( .D(n988), .CP(clk), .Q(\memory[19][35] ) );
  CFD1QXL \memory_reg[19][34]  ( .D(n989), .CP(clk), .Q(\memory[19][34] ) );
  CFD1QXL \memory_reg[19][33]  ( .D(n990), .CP(clk), .Q(\memory[19][33] ) );
  CFD1QXL \memory_reg[19][32]  ( .D(n991), .CP(clk), .Q(\memory[19][32] ) );
  CFD1QXL \memory_reg[19][31]  ( .D(n992), .CP(clk), .Q(\memory[19][31] ) );
  CFD1QXL \memory_reg[19][30]  ( .D(n993), .CP(clk), .Q(\memory[19][30] ) );
  CFD1QXL \memory_reg[19][29]  ( .D(n994), .CP(clk), .Q(\memory[19][29] ) );
  CFD1QXL \memory_reg[19][28]  ( .D(n995), .CP(clk), .Q(\memory[19][28] ) );
  CFD1QXL \memory_reg[19][27]  ( .D(n996), .CP(clk), .Q(\memory[19][27] ) );
  CFD1QXL \memory_reg[19][26]  ( .D(n997), .CP(clk), .Q(\memory[19][26] ) );
  CFD1QXL \memory_reg[19][25]  ( .D(n998), .CP(clk), .Q(\memory[19][25] ) );
  CFD1QXL \memory_reg[19][24]  ( .D(n999), .CP(clk), .Q(\memory[19][24] ) );
  CFD1QXL \memory_reg[19][23]  ( .D(n1000), .CP(clk), .Q(\memory[19][23] ) );
  CFD1QXL \memory_reg[19][22]  ( .D(n1001), .CP(clk), .Q(\memory[19][22] ) );
  CFD1QXL \memory_reg[19][21]  ( .D(n1002), .CP(clk), .Q(\memory[19][21] ) );
  CFD1QXL \memory_reg[19][20]  ( .D(n1003), .CP(clk), .Q(\memory[19][20] ) );
  CFD1QXL \memory_reg[19][19]  ( .D(n1004), .CP(clk), .Q(\memory[19][19] ) );
  CFD1QXL \memory_reg[19][18]  ( .D(n1005), .CP(clk), .Q(\memory[19][18] ) );
  CFD1QXL \memory_reg[19][17]  ( .D(n1006), .CP(clk), .Q(\memory[19][17] ) );
  CFD1QXL \memory_reg[19][16]  ( .D(n1007), .CP(clk), .Q(\memory[19][16] ) );
  CFD1QXL \memory_reg[19][15]  ( .D(n1008), .CP(clk), .Q(\memory[19][15] ) );
  CFD1QXL \memory_reg[19][14]  ( .D(n1009), .CP(clk), .Q(\memory[19][14] ) );
  CFD1QXL \memory_reg[19][13]  ( .D(n1010), .CP(clk), .Q(\memory[19][13] ) );
  CFD1QXL \memory_reg[19][12]  ( .D(n1011), .CP(clk), .Q(\memory[19][12] ) );
  CFD1QXL \memory_reg[19][11]  ( .D(n1012), .CP(clk), .Q(\memory[19][11] ) );
  CFD1QXL \memory_reg[19][10]  ( .D(n1013), .CP(clk), .Q(\memory[19][10] ) );
  CFD1QXL \memory_reg[19][9]  ( .D(n1014), .CP(clk), .Q(\memory[19][9] ) );
  CFD1QXL \memory_reg[19][8]  ( .D(n1015), .CP(clk), .Q(\memory[19][8] ) );
  CFD1QXL \memory_reg[19][7]  ( .D(n1016), .CP(clk), .Q(\memory[19][7] ) );
  CFD1QXL \memory_reg[19][6]  ( .D(n1017), .CP(clk), .Q(\memory[19][6] ) );
  CFD1QXL \memory_reg[19][5]  ( .D(n1018), .CP(clk), .Q(\memory[19][5] ) );
  CFD1QXL \memory_reg[19][4]  ( .D(n1019), .CP(clk), .Q(\memory[19][4] ) );
  CFD1QXL \memory_reg[19][3]  ( .D(n1020), .CP(clk), .Q(\memory[19][3] ) );
  CFD1QXL \memory_reg[19][2]  ( .D(n1021), .CP(clk), .Q(\memory[19][2] ) );
  CFD1QXL \memory_reg[19][1]  ( .D(n1022), .CP(clk), .Q(\memory[19][1] ) );
  CFD1QXL \memory_reg[19][0]  ( .D(n1023), .CP(clk), .Q(\memory[19][0] ) );
  CFD1QXL \memory_reg[15][63]  ( .D(n1244), .CP(clk), .Q(\memory[15][63] ) );
  CFD1QXL \memory_reg[15][61]  ( .D(n1246), .CP(clk), .Q(\memory[15][61] ) );
  CFD1QXL \memory_reg[15][60]  ( .D(n1247), .CP(clk), .Q(\memory[15][60] ) );
  CFD1QXL \memory_reg[15][59]  ( .D(n1248), .CP(clk), .Q(\memory[15][59] ) );
  CFD1QXL \memory_reg[15][58]  ( .D(n1249), .CP(clk), .Q(\memory[15][58] ) );
  CFD1QXL \memory_reg[15][57]  ( .D(n1250), .CP(clk), .Q(\memory[15][57] ) );
  CFD1QXL \memory_reg[15][56]  ( .D(n1251), .CP(clk), .Q(\memory[15][56] ) );
  CFD1QXL \memory_reg[15][55]  ( .D(n1252), .CP(clk), .Q(\memory[15][55] ) );
  CFD1QXL \memory_reg[15][54]  ( .D(n1253), .CP(clk), .Q(\memory[15][54] ) );
  CFD1QXL \memory_reg[15][53]  ( .D(n1254), .CP(clk), .Q(\memory[15][53] ) );
  CFD1QXL \memory_reg[15][52]  ( .D(n1255), .CP(clk), .Q(\memory[15][52] ) );
  CFD1QXL \memory_reg[15][51]  ( .D(n1256), .CP(clk), .Q(\memory[15][51] ) );
  CFD1QXL \memory_reg[15][50]  ( .D(n1257), .CP(clk), .Q(\memory[15][50] ) );
  CFD1QXL \memory_reg[15][49]  ( .D(n1258), .CP(clk), .Q(\memory[15][49] ) );
  CFD1QXL \memory_reg[15][48]  ( .D(n1259), .CP(clk), .Q(\memory[15][48] ) );
  CFD1QXL \memory_reg[15][47]  ( .D(n1260), .CP(clk), .Q(\memory[15][47] ) );
  CFD1QXL \memory_reg[15][46]  ( .D(n1261), .CP(clk), .Q(\memory[15][46] ) );
  CFD1QXL \memory_reg[15][45]  ( .D(n1262), .CP(clk), .Q(\memory[15][45] ) );
  CFD1QXL \memory_reg[15][44]  ( .D(n1263), .CP(clk), .Q(\memory[15][44] ) );
  CFD1QXL \memory_reg[15][43]  ( .D(n1264), .CP(clk), .Q(\memory[15][43] ) );
  CFD1QXL \memory_reg[15][42]  ( .D(n1265), .CP(clk), .Q(\memory[15][42] ) );
  CFD1QXL \memory_reg[15][41]  ( .D(n1266), .CP(clk), .Q(\memory[15][41] ) );
  CFD1QXL \memory_reg[15][40]  ( .D(n1267), .CP(clk), .Q(\memory[15][40] ) );
  CFD1QXL \memory_reg[15][39]  ( .D(n1268), .CP(clk), .Q(\memory[15][39] ) );
  CFD1QXL \memory_reg[15][38]  ( .D(n1269), .CP(clk), .Q(\memory[15][38] ) );
  CFD1QXL \memory_reg[15][37]  ( .D(n1270), .CP(clk), .Q(\memory[15][37] ) );
  CFD1QXL \memory_reg[15][36]  ( .D(n1271), .CP(clk), .Q(\memory[15][36] ) );
  CFD1QXL \memory_reg[15][35]  ( .D(n1272), .CP(clk), .Q(\memory[15][35] ) );
  CFD1QXL \memory_reg[15][34]  ( .D(n1273), .CP(clk), .Q(\memory[15][34] ) );
  CFD1QXL \memory_reg[15][33]  ( .D(n1274), .CP(clk), .Q(\memory[15][33] ) );
  CFD1QXL \memory_reg[15][32]  ( .D(n1275), .CP(clk), .Q(\memory[15][32] ) );
  CFD1QXL \memory_reg[15][31]  ( .D(n1276), .CP(clk), .Q(\memory[15][31] ) );
  CFD1QXL \memory_reg[15][30]  ( .D(n1277), .CP(clk), .Q(\memory[15][30] ) );
  CFD1QXL \memory_reg[15][29]  ( .D(n1278), .CP(clk), .Q(\memory[15][29] ) );
  CFD1QXL \memory_reg[15][28]  ( .D(n1279), .CP(clk), .Q(\memory[15][28] ) );
  CFD1QXL \memory_reg[15][27]  ( .D(n1280), .CP(clk), .Q(\memory[15][27] ) );
  CFD1QXL \memory_reg[15][26]  ( .D(n1281), .CP(clk), .Q(\memory[15][26] ) );
  CFD1QXL \memory_reg[15][25]  ( .D(n1282), .CP(clk), .Q(\memory[15][25] ) );
  CFD1QXL \memory_reg[15][24]  ( .D(n1283), .CP(clk), .Q(\memory[15][24] ) );
  CFD1QXL \memory_reg[15][23]  ( .D(n1284), .CP(clk), .Q(\memory[15][23] ) );
  CFD1QXL \memory_reg[15][22]  ( .D(n1285), .CP(clk), .Q(\memory[15][22] ) );
  CFD1QXL \memory_reg[15][21]  ( .D(n1286), .CP(clk), .Q(\memory[15][21] ) );
  CFD1QXL \memory_reg[15][20]  ( .D(n1287), .CP(clk), .Q(\memory[15][20] ) );
  CFD1QXL \memory_reg[15][19]  ( .D(n1288), .CP(clk), .Q(\memory[15][19] ) );
  CFD1QXL \memory_reg[15][18]  ( .D(n1289), .CP(clk), .Q(\memory[15][18] ) );
  CFD1QXL \memory_reg[15][17]  ( .D(n1290), .CP(clk), .Q(\memory[15][17] ) );
  CFD1QXL \memory_reg[15][16]  ( .D(n1291), .CP(clk), .Q(\memory[15][16] ) );
  CFD1QXL \memory_reg[15][15]  ( .D(n1292), .CP(clk), .Q(\memory[15][15] ) );
  CFD1QXL \memory_reg[15][14]  ( .D(n1293), .CP(clk), .Q(\memory[15][14] ) );
  CFD1QXL \memory_reg[15][13]  ( .D(n1294), .CP(clk), .Q(\memory[15][13] ) );
  CFD1QXL \memory_reg[15][12]  ( .D(n1295), .CP(clk), .Q(\memory[15][12] ) );
  CFD1QXL \memory_reg[15][11]  ( .D(n1296), .CP(clk), .Q(\memory[15][11] ) );
  CFD1QXL \memory_reg[15][10]  ( .D(n1297), .CP(clk), .Q(\memory[15][10] ) );
  CFD1QXL \memory_reg[15][9]  ( .D(n1298), .CP(clk), .Q(\memory[15][9] ) );
  CFD1QXL \memory_reg[15][8]  ( .D(n1299), .CP(clk), .Q(\memory[15][8] ) );
  CFD1QXL \memory_reg[15][7]  ( .D(n1300), .CP(clk), .Q(\memory[15][7] ) );
  CFD1QXL \memory_reg[15][6]  ( .D(n1301), .CP(clk), .Q(\memory[15][6] ) );
  CFD1QXL \memory_reg[15][5]  ( .D(n1302), .CP(clk), .Q(\memory[15][5] ) );
  CFD1QXL \memory_reg[15][4]  ( .D(n1303), .CP(clk), .Q(\memory[15][4] ) );
  CFD1QXL \memory_reg[15][3]  ( .D(n1304), .CP(clk), .Q(\memory[15][3] ) );
  CFD1QXL \memory_reg[15][2]  ( .D(n1305), .CP(clk), .Q(\memory[15][2] ) );
  CFD1QXL \memory_reg[15][1]  ( .D(n1306), .CP(clk), .Q(\memory[15][1] ) );
  CFD1QXL \memory_reg[15][0]  ( .D(n1307), .CP(clk), .Q(\memory[15][0] ) );
  CFD1QXL \memory_reg[30][63]  ( .D(n179), .CP(clk), .Q(\memory[30][63] ) );
  CFD1QXL \memory_reg[30][62]  ( .D(n180), .CP(clk), .Q(\memory[30][62] ) );
  CFD1QXL \memory_reg[30][61]  ( .D(n181), .CP(clk), .Q(\memory[30][61] ) );
  CFD1QXL \memory_reg[30][60]  ( .D(n182), .CP(clk), .Q(\memory[30][60] ) );
  CFD1QXL \memory_reg[30][59]  ( .D(n183), .CP(clk), .Q(\memory[30][59] ) );
  CFD1QXL \memory_reg[30][58]  ( .D(n184), .CP(clk), .Q(\memory[30][58] ) );
  CFD1QXL \memory_reg[30][57]  ( .D(n185), .CP(clk), .Q(\memory[30][57] ) );
  CFD1QXL \memory_reg[30][56]  ( .D(n186), .CP(clk), .Q(\memory[30][56] ) );
  CFD1QXL \memory_reg[30][55]  ( .D(n187), .CP(clk), .Q(\memory[30][55] ) );
  CFD1QXL \memory_reg[30][54]  ( .D(n188), .CP(clk), .Q(\memory[30][54] ) );
  CFD1QXL \memory_reg[30][53]  ( .D(n189), .CP(clk), .Q(\memory[30][53] ) );
  CFD1QXL \memory_reg[30][52]  ( .D(n190), .CP(clk), .Q(\memory[30][52] ) );
  CFD1QXL \memory_reg[30][51]  ( .D(n191), .CP(clk), .Q(\memory[30][51] ) );
  CFD1QXL \memory_reg[30][50]  ( .D(n192), .CP(clk), .Q(\memory[30][50] ) );
  CFD1QXL \memory_reg[30][49]  ( .D(n193), .CP(clk), .Q(\memory[30][49] ) );
  CFD1QXL \memory_reg[30][48]  ( .D(n194), .CP(clk), .Q(\memory[30][48] ) );
  CFD1QXL \memory_reg[30][47]  ( .D(n195), .CP(clk), .Q(\memory[30][47] ) );
  CFD1QXL \memory_reg[30][46]  ( .D(n196), .CP(clk), .Q(\memory[30][46] ) );
  CFD1QXL \memory_reg[30][45]  ( .D(n197), .CP(clk), .Q(\memory[30][45] ) );
  CFD1QXL \memory_reg[30][44]  ( .D(n198), .CP(clk), .Q(\memory[30][44] ) );
  CFD1QXL \memory_reg[30][43]  ( .D(n199), .CP(clk), .Q(\memory[30][43] ) );
  CFD1QXL \memory_reg[30][42]  ( .D(n200), .CP(clk), .Q(\memory[30][42] ) );
  CFD1QXL \memory_reg[30][41]  ( .D(n201), .CP(clk), .Q(\memory[30][41] ) );
  CFD1QXL \memory_reg[30][40]  ( .D(n202), .CP(clk), .Q(\memory[30][40] ) );
  CFD1QXL \memory_reg[30][39]  ( .D(n203), .CP(clk), .Q(\memory[30][39] ) );
  CFD1QXL \memory_reg[30][38]  ( .D(n204), .CP(clk), .Q(\memory[30][38] ) );
  CFD1QXL \memory_reg[30][37]  ( .D(n205), .CP(clk), .Q(\memory[30][37] ) );
  CFD1QXL \memory_reg[30][36]  ( .D(n206), .CP(clk), .Q(\memory[30][36] ) );
  CFD1QXL \memory_reg[30][35]  ( .D(n207), .CP(clk), .Q(\memory[30][35] ) );
  CFD1QXL \memory_reg[30][34]  ( .D(n208), .CP(clk), .Q(\memory[30][34] ) );
  CFD1QXL \memory_reg[30][33]  ( .D(n209), .CP(clk), .Q(\memory[30][33] ) );
  CFD1QXL \memory_reg[30][32]  ( .D(n210), .CP(clk), .Q(\memory[30][32] ) );
  CFD1QXL \memory_reg[30][31]  ( .D(n211), .CP(clk), .Q(\memory[30][31] ) );
  CFD1QXL \memory_reg[30][30]  ( .D(n212), .CP(clk), .Q(\memory[30][30] ) );
  CFD1QXL \memory_reg[30][29]  ( .D(n213), .CP(clk), .Q(\memory[30][29] ) );
  CFD1QXL \memory_reg[30][28]  ( .D(n214), .CP(clk), .Q(\memory[30][28] ) );
  CFD1QXL \memory_reg[30][27]  ( .D(n215), .CP(clk), .Q(\memory[30][27] ) );
  CFD1QXL \memory_reg[30][26]  ( .D(n216), .CP(clk), .Q(\memory[30][26] ) );
  CFD1QXL \memory_reg[30][25]  ( .D(n217), .CP(clk), .Q(\memory[30][25] ) );
  CFD1QXL \memory_reg[30][24]  ( .D(n218), .CP(clk), .Q(\memory[30][24] ) );
  CFD1QXL \memory_reg[30][23]  ( .D(n219), .CP(clk), .Q(\memory[30][23] ) );
  CFD1QXL \memory_reg[30][22]  ( .D(n220), .CP(clk), .Q(\memory[30][22] ) );
  CFD1QXL \memory_reg[30][21]  ( .D(n221), .CP(clk), .Q(\memory[30][21] ) );
  CFD1QXL \memory_reg[30][20]  ( .D(n222), .CP(clk), .Q(\memory[30][20] ) );
  CFD1QXL \memory_reg[30][19]  ( .D(n223), .CP(clk), .Q(\memory[30][19] ) );
  CFD1QXL \memory_reg[30][18]  ( .D(n224), .CP(clk), .Q(\memory[30][18] ) );
  CFD1QXL \memory_reg[30][17]  ( .D(n225), .CP(clk), .Q(\memory[30][17] ) );
  CFD1QXL \memory_reg[30][16]  ( .D(n226), .CP(clk), .Q(\memory[30][16] ) );
  CFD1QXL \memory_reg[30][15]  ( .D(n227), .CP(clk), .Q(\memory[30][15] ) );
  CFD1QXL \memory_reg[30][14]  ( .D(n228), .CP(clk), .Q(\memory[30][14] ) );
  CFD1QXL \memory_reg[30][13]  ( .D(n229), .CP(clk), .Q(\memory[30][13] ) );
  CFD1QXL \memory_reg[30][12]  ( .D(n230), .CP(clk), .Q(\memory[30][12] ) );
  CFD1QXL \memory_reg[30][11]  ( .D(n231), .CP(clk), .Q(\memory[30][11] ) );
  CFD1QXL \memory_reg[30][10]  ( .D(n232), .CP(clk), .Q(\memory[30][10] ) );
  CFD1QXL \memory_reg[30][9]  ( .D(n233), .CP(clk), .Q(\memory[30][9] ) );
  CFD1QXL \memory_reg[30][8]  ( .D(n234), .CP(clk), .Q(\memory[30][8] ) );
  CFD1QXL \memory_reg[30][7]  ( .D(n235), .CP(clk), .Q(\memory[30][7] ) );
  CFD1QXL \memory_reg[30][6]  ( .D(n236), .CP(clk), .Q(\memory[30][6] ) );
  CFD1QXL \memory_reg[30][5]  ( .D(n237), .CP(clk), .Q(\memory[30][5] ) );
  CFD1QXL \memory_reg[30][4]  ( .D(n238), .CP(clk), .Q(\memory[30][4] ) );
  CFD1QXL \memory_reg[30][3]  ( .D(n239), .CP(clk), .Q(\memory[30][3] ) );
  CFD1QXL \memory_reg[30][2]  ( .D(n240), .CP(clk), .Q(\memory[30][2] ) );
  CFD1QXL \memory_reg[30][1]  ( .D(n241), .CP(clk), .Q(\memory[30][1] ) );
  CFD1QXL \memory_reg[30][0]  ( .D(n242), .CP(clk), .Q(\memory[30][0] ) );
  CFD1QXL \memory_reg[29][63]  ( .D(n250), .CP(clk), .Q(\memory[29][63] ) );
  CFD1QXL \memory_reg[29][62]  ( .D(n251), .CP(clk), .Q(\memory[29][62] ) );
  CFD1QXL \memory_reg[29][61]  ( .D(n252), .CP(clk), .Q(\memory[29][61] ) );
  CFD1QXL \memory_reg[29][60]  ( .D(n253), .CP(clk), .Q(\memory[29][60] ) );
  CFD1QXL \memory_reg[29][59]  ( .D(n254), .CP(clk), .Q(\memory[29][59] ) );
  CFD1QXL \memory_reg[29][58]  ( .D(n255), .CP(clk), .Q(\memory[29][58] ) );
  CFD1QXL \memory_reg[29][57]  ( .D(n256), .CP(clk), .Q(\memory[29][57] ) );
  CFD1QXL \memory_reg[29][56]  ( .D(n257), .CP(clk), .Q(\memory[29][56] ) );
  CFD1QXL \memory_reg[29][55]  ( .D(n258), .CP(clk), .Q(\memory[29][55] ) );
  CFD1QXL \memory_reg[29][54]  ( .D(n259), .CP(clk), .Q(\memory[29][54] ) );
  CFD1QXL \memory_reg[29][53]  ( .D(n260), .CP(clk), .Q(\memory[29][53] ) );
  CFD1QXL \memory_reg[29][52]  ( .D(n261), .CP(clk), .Q(\memory[29][52] ) );
  CFD1QXL \memory_reg[29][51]  ( .D(n262), .CP(clk), .Q(\memory[29][51] ) );
  CFD1QXL \memory_reg[29][50]  ( .D(n263), .CP(clk), .Q(\memory[29][50] ) );
  CFD1QXL \memory_reg[29][49]  ( .D(n264), .CP(clk), .Q(\memory[29][49] ) );
  CFD1QXL \memory_reg[29][48]  ( .D(n265), .CP(clk), .Q(\memory[29][48] ) );
  CFD1QXL \memory_reg[29][47]  ( .D(n266), .CP(clk), .Q(\memory[29][47] ) );
  CFD1QXL \memory_reg[29][46]  ( .D(n267), .CP(clk), .Q(\memory[29][46] ) );
  CFD1QXL \memory_reg[29][45]  ( .D(n268), .CP(clk), .Q(\memory[29][45] ) );
  CFD1QXL \memory_reg[29][44]  ( .D(n269), .CP(clk), .Q(\memory[29][44] ) );
  CFD1QXL \memory_reg[29][43]  ( .D(n270), .CP(clk), .Q(\memory[29][43] ) );
  CFD1QXL \memory_reg[29][42]  ( .D(n271), .CP(clk), .Q(\memory[29][42] ) );
  CFD1QXL \memory_reg[29][41]  ( .D(n272), .CP(clk), .Q(\memory[29][41] ) );
  CFD1QXL \memory_reg[29][40]  ( .D(n273), .CP(clk), .Q(\memory[29][40] ) );
  CFD1QXL \memory_reg[29][39]  ( .D(n274), .CP(clk), .Q(\memory[29][39] ) );
  CFD1QXL \memory_reg[29][38]  ( .D(n275), .CP(clk), .Q(\memory[29][38] ) );
  CFD1QXL \memory_reg[29][37]  ( .D(n276), .CP(clk), .Q(\memory[29][37] ) );
  CFD1QXL \memory_reg[29][36]  ( .D(n277), .CP(clk), .Q(\memory[29][36] ) );
  CFD1QXL \memory_reg[29][35]  ( .D(n278), .CP(clk), .Q(\memory[29][35] ) );
  CFD1QXL \memory_reg[29][34]  ( .D(n279), .CP(clk), .Q(\memory[29][34] ) );
  CFD1QXL \memory_reg[29][33]  ( .D(n280), .CP(clk), .Q(\memory[29][33] ) );
  CFD1QXL \memory_reg[29][32]  ( .D(n281), .CP(clk), .Q(\memory[29][32] ) );
  CFD1QXL \memory_reg[29][31]  ( .D(n282), .CP(clk), .Q(\memory[29][31] ) );
  CFD1QXL \memory_reg[29][30]  ( .D(n283), .CP(clk), .Q(\memory[29][30] ) );
  CFD1QXL \memory_reg[29][29]  ( .D(n284), .CP(clk), .Q(\memory[29][29] ) );
  CFD1QXL \memory_reg[29][28]  ( .D(n285), .CP(clk), .Q(\memory[29][28] ) );
  CFD1QXL \memory_reg[29][27]  ( .D(n286), .CP(clk), .Q(\memory[29][27] ) );
  CFD1QXL \memory_reg[29][26]  ( .D(n287), .CP(clk), .Q(\memory[29][26] ) );
  CFD1QXL \memory_reg[29][25]  ( .D(n288), .CP(clk), .Q(\memory[29][25] ) );
  CFD1QXL \memory_reg[29][24]  ( .D(n289), .CP(clk), .Q(\memory[29][24] ) );
  CFD1QXL \memory_reg[29][23]  ( .D(n290), .CP(clk), .Q(\memory[29][23] ) );
  CFD1QXL \memory_reg[29][22]  ( .D(n291), .CP(clk), .Q(\memory[29][22] ) );
  CFD1QXL \memory_reg[29][21]  ( .D(n292), .CP(clk), .Q(\memory[29][21] ) );
  CFD1QXL \memory_reg[29][20]  ( .D(n293), .CP(clk), .Q(\memory[29][20] ) );
  CFD1QXL \memory_reg[29][19]  ( .D(n294), .CP(clk), .Q(\memory[29][19] ) );
  CFD1QXL \memory_reg[29][18]  ( .D(n295), .CP(clk), .Q(\memory[29][18] ) );
  CFD1QXL \memory_reg[29][17]  ( .D(n296), .CP(clk), .Q(\memory[29][17] ) );
  CFD1QXL \memory_reg[29][16]  ( .D(n297), .CP(clk), .Q(\memory[29][16] ) );
  CFD1QXL \memory_reg[29][15]  ( .D(n298), .CP(clk), .Q(\memory[29][15] ) );
  CFD1QXL \memory_reg[29][14]  ( .D(n299), .CP(clk), .Q(\memory[29][14] ) );
  CFD1QXL \memory_reg[29][13]  ( .D(n300), .CP(clk), .Q(\memory[29][13] ) );
  CFD1QXL \memory_reg[29][12]  ( .D(n301), .CP(clk), .Q(\memory[29][12] ) );
  CFD1QXL \memory_reg[29][11]  ( .D(n302), .CP(clk), .Q(\memory[29][11] ) );
  CFD1QXL \memory_reg[29][10]  ( .D(n303), .CP(clk), .Q(\memory[29][10] ) );
  CFD1QXL \memory_reg[29][9]  ( .D(n304), .CP(clk), .Q(\memory[29][9] ) );
  CFD1QXL \memory_reg[29][8]  ( .D(n305), .CP(clk), .Q(\memory[29][8] ) );
  CFD1QXL \memory_reg[29][7]  ( .D(n306), .CP(clk), .Q(\memory[29][7] ) );
  CFD1QXL \memory_reg[29][6]  ( .D(n307), .CP(clk), .Q(\memory[29][6] ) );
  CFD1QXL \memory_reg[29][5]  ( .D(n308), .CP(clk), .Q(\memory[29][5] ) );
  CFD1QXL \memory_reg[29][4]  ( .D(n309), .CP(clk), .Q(\memory[29][4] ) );
  CFD1QXL \memory_reg[29][3]  ( .D(n310), .CP(clk), .Q(\memory[29][3] ) );
  CFD1QXL \memory_reg[29][2]  ( .D(n311), .CP(clk), .Q(\memory[29][2] ) );
  CFD1QXL \memory_reg[29][1]  ( .D(n312), .CP(clk), .Q(\memory[29][1] ) );
  CFD1QXL \memory_reg[29][0]  ( .D(n313), .CP(clk), .Q(\memory[29][0] ) );
  CFD1QXL \memory_reg[28][63]  ( .D(n321), .CP(clk), .Q(\memory[28][63] ) );
  CFD1QXL \memory_reg[28][62]  ( .D(n322), .CP(clk), .Q(\memory[28][62] ) );
  CFD1QXL \memory_reg[28][61]  ( .D(n323), .CP(clk), .Q(\memory[28][61] ) );
  CFD1QXL \memory_reg[28][60]  ( .D(n324), .CP(clk), .Q(\memory[28][60] ) );
  CFD1QXL \memory_reg[28][59]  ( .D(n325), .CP(clk), .Q(\memory[28][59] ) );
  CFD1QXL \memory_reg[28][58]  ( .D(n326), .CP(clk), .Q(\memory[28][58] ) );
  CFD1QXL \memory_reg[28][57]  ( .D(n327), .CP(clk), .Q(\memory[28][57] ) );
  CFD1QXL \memory_reg[28][56]  ( .D(n328), .CP(clk), .Q(\memory[28][56] ) );
  CFD1QXL \memory_reg[28][55]  ( .D(n329), .CP(clk), .Q(\memory[28][55] ) );
  CFD1QXL \memory_reg[28][54]  ( .D(n330), .CP(clk), .Q(\memory[28][54] ) );
  CFD1QXL \memory_reg[28][53]  ( .D(n331), .CP(clk), .Q(\memory[28][53] ) );
  CFD1QXL \memory_reg[28][52]  ( .D(n332), .CP(clk), .Q(\memory[28][52] ) );
  CFD1QXL \memory_reg[28][51]  ( .D(n333), .CP(clk), .Q(\memory[28][51] ) );
  CFD1QXL \memory_reg[28][50]  ( .D(n334), .CP(clk), .Q(\memory[28][50] ) );
  CFD1QXL \memory_reg[28][49]  ( .D(n335), .CP(clk), .Q(\memory[28][49] ) );
  CFD1QXL \memory_reg[28][48]  ( .D(n336), .CP(clk), .Q(\memory[28][48] ) );
  CFD1QXL \memory_reg[28][47]  ( .D(n337), .CP(clk), .Q(\memory[28][47] ) );
  CFD1QXL \memory_reg[28][46]  ( .D(n338), .CP(clk), .Q(\memory[28][46] ) );
  CFD1QXL \memory_reg[28][45]  ( .D(n339), .CP(clk), .Q(\memory[28][45] ) );
  CFD1QXL \memory_reg[28][44]  ( .D(n340), .CP(clk), .Q(\memory[28][44] ) );
  CFD1QXL \memory_reg[28][43]  ( .D(n341), .CP(clk), .Q(\memory[28][43] ) );
  CFD1QXL \memory_reg[28][42]  ( .D(n342), .CP(clk), .Q(\memory[28][42] ) );
  CFD1QXL \memory_reg[28][41]  ( .D(n343), .CP(clk), .Q(\memory[28][41] ) );
  CFD1QXL \memory_reg[28][40]  ( .D(n344), .CP(clk), .Q(\memory[28][40] ) );
  CFD1QXL \memory_reg[28][39]  ( .D(n345), .CP(clk), .Q(\memory[28][39] ) );
  CFD1QXL \memory_reg[28][38]  ( .D(n346), .CP(clk), .Q(\memory[28][38] ) );
  CFD1QXL \memory_reg[28][37]  ( .D(n347), .CP(clk), .Q(\memory[28][37] ) );
  CFD1QXL \memory_reg[28][36]  ( .D(n348), .CP(clk), .Q(\memory[28][36] ) );
  CFD1QXL \memory_reg[28][35]  ( .D(n349), .CP(clk), .Q(\memory[28][35] ) );
  CFD1QXL \memory_reg[28][34]  ( .D(n350), .CP(clk), .Q(\memory[28][34] ) );
  CFD1QXL \memory_reg[28][33]  ( .D(n351), .CP(clk), .Q(\memory[28][33] ) );
  CFD1QXL \memory_reg[28][32]  ( .D(n352), .CP(clk), .Q(\memory[28][32] ) );
  CFD1QXL \memory_reg[28][31]  ( .D(n353), .CP(clk), .Q(\memory[28][31] ) );
  CFD1QXL \memory_reg[28][30]  ( .D(n354), .CP(clk), .Q(\memory[28][30] ) );
  CFD1QXL \memory_reg[28][29]  ( .D(n355), .CP(clk), .Q(\memory[28][29] ) );
  CFD1QXL \memory_reg[28][28]  ( .D(n356), .CP(clk), .Q(\memory[28][28] ) );
  CFD1QXL \memory_reg[28][27]  ( .D(n357), .CP(clk), .Q(\memory[28][27] ) );
  CFD1QXL \memory_reg[28][26]  ( .D(n358), .CP(clk), .Q(\memory[28][26] ) );
  CFD1QXL \memory_reg[28][25]  ( .D(n359), .CP(clk), .Q(\memory[28][25] ) );
  CFD1QXL \memory_reg[28][24]  ( .D(n360), .CP(clk), .Q(\memory[28][24] ) );
  CFD1QXL \memory_reg[28][23]  ( .D(n361), .CP(clk), .Q(\memory[28][23] ) );
  CFD1QXL \memory_reg[28][22]  ( .D(n362), .CP(clk), .Q(\memory[28][22] ) );
  CFD1QXL \memory_reg[28][21]  ( .D(n363), .CP(clk), .Q(\memory[28][21] ) );
  CFD1QXL \memory_reg[28][20]  ( .D(n364), .CP(clk), .Q(\memory[28][20] ) );
  CFD1QXL \memory_reg[28][19]  ( .D(n365), .CP(clk), .Q(\memory[28][19] ) );
  CFD1QXL \memory_reg[28][18]  ( .D(n366), .CP(clk), .Q(\memory[28][18] ) );
  CFD1QXL \memory_reg[28][17]  ( .D(n367), .CP(clk), .Q(\memory[28][17] ) );
  CFD1QXL \memory_reg[28][16]  ( .D(n368), .CP(clk), .Q(\memory[28][16] ) );
  CFD1QXL \memory_reg[28][15]  ( .D(n369), .CP(clk), .Q(\memory[28][15] ) );
  CFD1QXL \memory_reg[28][14]  ( .D(n370), .CP(clk), .Q(\memory[28][14] ) );
  CFD1QXL \memory_reg[28][13]  ( .D(n371), .CP(clk), .Q(\memory[28][13] ) );
  CFD1QXL \memory_reg[28][12]  ( .D(n372), .CP(clk), .Q(\memory[28][12] ) );
  CFD1QXL \memory_reg[28][11]  ( .D(n373), .CP(clk), .Q(\memory[28][11] ) );
  CFD1QXL \memory_reg[28][10]  ( .D(n374), .CP(clk), .Q(\memory[28][10] ) );
  CFD1QXL \memory_reg[28][9]  ( .D(n375), .CP(clk), .Q(\memory[28][9] ) );
  CFD1QXL \memory_reg[28][8]  ( .D(n376), .CP(clk), .Q(\memory[28][8] ) );
  CFD1QXL \memory_reg[28][7]  ( .D(n377), .CP(clk), .Q(\memory[28][7] ) );
  CFD1QXL \memory_reg[28][6]  ( .D(n378), .CP(clk), .Q(\memory[28][6] ) );
  CFD1QXL \memory_reg[28][5]  ( .D(n379), .CP(clk), .Q(\memory[28][5] ) );
  CFD1QXL \memory_reg[28][4]  ( .D(n380), .CP(clk), .Q(\memory[28][4] ) );
  CFD1QXL \memory_reg[28][3]  ( .D(n381), .CP(clk), .Q(\memory[28][3] ) );
  CFD1QXL \memory_reg[28][2]  ( .D(n382), .CP(clk), .Q(\memory[28][2] ) );
  CFD1QXL \memory_reg[28][1]  ( .D(n383), .CP(clk), .Q(\memory[28][1] ) );
  CFD1QXL \memory_reg[28][0]  ( .D(n384), .CP(clk), .Q(\memory[28][0] ) );
  CFD1QXL \memory_reg[26][63]  ( .D(n463), .CP(clk), .Q(\memory[26][63] ) );
  CFD1QXL \memory_reg[26][62]  ( .D(n464), .CP(clk), .Q(\memory[26][62] ) );
  CFD1QXL \memory_reg[26][61]  ( .D(n465), .CP(clk), .Q(\memory[26][61] ) );
  CFD1QXL \memory_reg[26][60]  ( .D(n466), .CP(clk), .Q(\memory[26][60] ) );
  CFD1QXL \memory_reg[26][59]  ( .D(n467), .CP(clk), .Q(\memory[26][59] ) );
  CFD1QXL \memory_reg[26][58]  ( .D(n468), .CP(clk), .Q(\memory[26][58] ) );
  CFD1QXL \memory_reg[26][57]  ( .D(n469), .CP(clk), .Q(\memory[26][57] ) );
  CFD1QXL \memory_reg[26][56]  ( .D(n470), .CP(clk), .Q(\memory[26][56] ) );
  CFD1QXL \memory_reg[26][55]  ( .D(n471), .CP(clk), .Q(\memory[26][55] ) );
  CFD1QXL \memory_reg[26][54]  ( .D(n472), .CP(clk), .Q(\memory[26][54] ) );
  CFD1QXL \memory_reg[26][53]  ( .D(n473), .CP(clk), .Q(\memory[26][53] ) );
  CFD1QXL \memory_reg[26][52]  ( .D(n474), .CP(clk), .Q(\memory[26][52] ) );
  CFD1QXL \memory_reg[26][51]  ( .D(n475), .CP(clk), .Q(\memory[26][51] ) );
  CFD1QXL \memory_reg[26][50]  ( .D(n476), .CP(clk), .Q(\memory[26][50] ) );
  CFD1QXL \memory_reg[26][49]  ( .D(n477), .CP(clk), .Q(\memory[26][49] ) );
  CFD1QXL \memory_reg[26][48]  ( .D(n478), .CP(clk), .Q(\memory[26][48] ) );
  CFD1QXL \memory_reg[26][47]  ( .D(n479), .CP(clk), .Q(\memory[26][47] ) );
  CFD1QXL \memory_reg[26][46]  ( .D(n480), .CP(clk), .Q(\memory[26][46] ) );
  CFD1QXL \memory_reg[26][45]  ( .D(n481), .CP(clk), .Q(\memory[26][45] ) );
  CFD1QXL \memory_reg[26][44]  ( .D(n482), .CP(clk), .Q(\memory[26][44] ) );
  CFD1QXL \memory_reg[26][43]  ( .D(n483), .CP(clk), .Q(\memory[26][43] ) );
  CFD1QXL \memory_reg[26][42]  ( .D(n484), .CP(clk), .Q(\memory[26][42] ) );
  CFD1QXL \memory_reg[26][41]  ( .D(n485), .CP(clk), .Q(\memory[26][41] ) );
  CFD1QXL \memory_reg[26][40]  ( .D(n486), .CP(clk), .Q(\memory[26][40] ) );
  CFD1QXL \memory_reg[26][39]  ( .D(n487), .CP(clk), .Q(\memory[26][39] ) );
  CFD1QXL \memory_reg[26][38]  ( .D(n488), .CP(clk), .Q(\memory[26][38] ) );
  CFD1QXL \memory_reg[26][37]  ( .D(n489), .CP(clk), .Q(\memory[26][37] ) );
  CFD1QXL \memory_reg[26][36]  ( .D(n490), .CP(clk), .Q(\memory[26][36] ) );
  CFD1QXL \memory_reg[26][35]  ( .D(n491), .CP(clk), .Q(\memory[26][35] ) );
  CFD1QXL \memory_reg[26][34]  ( .D(n492), .CP(clk), .Q(\memory[26][34] ) );
  CFD1QXL \memory_reg[26][33]  ( .D(n493), .CP(clk), .Q(\memory[26][33] ) );
  CFD1QXL \memory_reg[26][32]  ( .D(n494), .CP(clk), .Q(\memory[26][32] ) );
  CFD1QXL \memory_reg[26][31]  ( .D(n495), .CP(clk), .Q(\memory[26][31] ) );
  CFD1QXL \memory_reg[26][30]  ( .D(n496), .CP(clk), .Q(\memory[26][30] ) );
  CFD1QXL \memory_reg[26][29]  ( .D(n497), .CP(clk), .Q(\memory[26][29] ) );
  CFD1QXL \memory_reg[26][28]  ( .D(n498), .CP(clk), .Q(\memory[26][28] ) );
  CFD1QXL \memory_reg[26][27]  ( .D(n499), .CP(clk), .Q(\memory[26][27] ) );
  CFD1QXL \memory_reg[26][26]  ( .D(n500), .CP(clk), .Q(\memory[26][26] ) );
  CFD1QXL \memory_reg[26][25]  ( .D(n501), .CP(clk), .Q(\memory[26][25] ) );
  CFD1QXL \memory_reg[26][24]  ( .D(n502), .CP(clk), .Q(\memory[26][24] ) );
  CFD1QXL \memory_reg[26][23]  ( .D(n503), .CP(clk), .Q(\memory[26][23] ) );
  CFD1QXL \memory_reg[26][22]  ( .D(n504), .CP(clk), .Q(\memory[26][22] ) );
  CFD1QXL \memory_reg[26][21]  ( .D(n505), .CP(clk), .Q(\memory[26][21] ) );
  CFD1QXL \memory_reg[26][20]  ( .D(n506), .CP(clk), .Q(\memory[26][20] ) );
  CFD1QXL \memory_reg[26][19]  ( .D(n507), .CP(clk), .Q(\memory[26][19] ) );
  CFD1QXL \memory_reg[26][18]  ( .D(n508), .CP(clk), .Q(\memory[26][18] ) );
  CFD1QXL \memory_reg[26][17]  ( .D(n509), .CP(clk), .Q(\memory[26][17] ) );
  CFD1QXL \memory_reg[26][16]  ( .D(n510), .CP(clk), .Q(\memory[26][16] ) );
  CFD1QXL \memory_reg[26][15]  ( .D(n511), .CP(clk), .Q(\memory[26][15] ) );
  CFD1QXL \memory_reg[26][14]  ( .D(n512), .CP(clk), .Q(\memory[26][14] ) );
  CFD1QXL \memory_reg[26][13]  ( .D(n513), .CP(clk), .Q(\memory[26][13] ) );
  CFD1QXL \memory_reg[26][12]  ( .D(n514), .CP(clk), .Q(\memory[26][12] ) );
  CFD1QXL \memory_reg[26][11]  ( .D(n515), .CP(clk), .Q(\memory[26][11] ) );
  CFD1QXL \memory_reg[26][10]  ( .D(n516), .CP(clk), .Q(\memory[26][10] ) );
  CFD1QXL \memory_reg[26][9]  ( .D(n517), .CP(clk), .Q(\memory[26][9] ) );
  CFD1QXL \memory_reg[26][8]  ( .D(n518), .CP(clk), .Q(\memory[26][8] ) );
  CFD1QXL \memory_reg[26][7]  ( .D(n519), .CP(clk), .Q(\memory[26][7] ) );
  CFD1QXL \memory_reg[26][6]  ( .D(n520), .CP(clk), .Q(\memory[26][6] ) );
  CFD1QXL \memory_reg[26][5]  ( .D(n521), .CP(clk), .Q(\memory[26][5] ) );
  CFD1QXL \memory_reg[26][4]  ( .D(n522), .CP(clk), .Q(\memory[26][4] ) );
  CFD1QXL \memory_reg[26][3]  ( .D(n523), .CP(clk), .Q(\memory[26][3] ) );
  CFD1QXL \memory_reg[26][2]  ( .D(n524), .CP(clk), .Q(\memory[26][2] ) );
  CFD1QXL \memory_reg[26][1]  ( .D(n525), .CP(clk), .Q(\memory[26][1] ) );
  CFD1QXL \memory_reg[26][0]  ( .D(n526), .CP(clk), .Q(\memory[26][0] ) );
  CFD1QXL \memory_reg[25][63]  ( .D(n534), .CP(clk), .Q(\memory[25][63] ) );
  CFD1QXL \memory_reg[25][62]  ( .D(n535), .CP(clk), .Q(\memory[25][62] ) );
  CFD1QXL \memory_reg[25][61]  ( .D(n536), .CP(clk), .Q(\memory[25][61] ) );
  CFD1QXL \memory_reg[25][60]  ( .D(n537), .CP(clk), .Q(\memory[25][60] ) );
  CFD1QXL \memory_reg[25][59]  ( .D(n538), .CP(clk), .Q(\memory[25][59] ) );
  CFD1QXL \memory_reg[25][58]  ( .D(n539), .CP(clk), .Q(\memory[25][58] ) );
  CFD1QXL \memory_reg[25][57]  ( .D(n540), .CP(clk), .Q(\memory[25][57] ) );
  CFD1QXL \memory_reg[25][56]  ( .D(n541), .CP(clk), .Q(\memory[25][56] ) );
  CFD1QXL \memory_reg[25][55]  ( .D(n542), .CP(clk), .Q(\memory[25][55] ) );
  CFD1QXL \memory_reg[25][54]  ( .D(n543), .CP(clk), .Q(\memory[25][54] ) );
  CFD1QXL \memory_reg[25][53]  ( .D(n544), .CP(clk), .Q(\memory[25][53] ) );
  CFD1QXL \memory_reg[25][52]  ( .D(n545), .CP(clk), .Q(\memory[25][52] ) );
  CFD1QXL \memory_reg[25][51]  ( .D(n546), .CP(clk), .Q(\memory[25][51] ) );
  CFD1QXL \memory_reg[25][50]  ( .D(n547), .CP(clk), .Q(\memory[25][50] ) );
  CFD1QXL \memory_reg[25][49]  ( .D(n548), .CP(clk), .Q(\memory[25][49] ) );
  CFD1QXL \memory_reg[25][48]  ( .D(n549), .CP(clk), .Q(\memory[25][48] ) );
  CFD1QXL \memory_reg[25][47]  ( .D(n550), .CP(clk), .Q(\memory[25][47] ) );
  CFD1QXL \memory_reg[25][46]  ( .D(n551), .CP(clk), .Q(\memory[25][46] ) );
  CFD1QXL \memory_reg[25][45]  ( .D(n552), .CP(clk), .Q(\memory[25][45] ) );
  CFD1QXL \memory_reg[25][44]  ( .D(n553), .CP(clk), .Q(\memory[25][44] ) );
  CFD1QXL \memory_reg[25][43]  ( .D(n554), .CP(clk), .Q(\memory[25][43] ) );
  CFD1QXL \memory_reg[25][42]  ( .D(n555), .CP(clk), .Q(\memory[25][42] ) );
  CFD1QXL \memory_reg[25][41]  ( .D(n556), .CP(clk), .Q(\memory[25][41] ) );
  CFD1QXL \memory_reg[25][40]  ( .D(n557), .CP(clk), .Q(\memory[25][40] ) );
  CFD1QXL \memory_reg[25][39]  ( .D(n558), .CP(clk), .Q(\memory[25][39] ) );
  CFD1QXL \memory_reg[25][38]  ( .D(n559), .CP(clk), .Q(\memory[25][38] ) );
  CFD1QXL \memory_reg[25][37]  ( .D(n560), .CP(clk), .Q(\memory[25][37] ) );
  CFD1QXL \memory_reg[25][36]  ( .D(n561), .CP(clk), .Q(\memory[25][36] ) );
  CFD1QXL \memory_reg[25][35]  ( .D(n562), .CP(clk), .Q(\memory[25][35] ) );
  CFD1QXL \memory_reg[25][34]  ( .D(n563), .CP(clk), .Q(\memory[25][34] ) );
  CFD1QXL \memory_reg[25][33]  ( .D(n564), .CP(clk), .Q(\memory[25][33] ) );
  CFD1QXL \memory_reg[25][32]  ( .D(n565), .CP(clk), .Q(\memory[25][32] ) );
  CFD1QXL \memory_reg[25][31]  ( .D(n566), .CP(clk), .Q(\memory[25][31] ) );
  CFD1QXL \memory_reg[25][30]  ( .D(n567), .CP(clk), .Q(\memory[25][30] ) );
  CFD1QXL \memory_reg[25][29]  ( .D(n568), .CP(clk), .Q(\memory[25][29] ) );
  CFD1QXL \memory_reg[25][28]  ( .D(n569), .CP(clk), .Q(\memory[25][28] ) );
  CFD1QXL \memory_reg[25][27]  ( .D(n570), .CP(clk), .Q(\memory[25][27] ) );
  CFD1QXL \memory_reg[25][26]  ( .D(n571), .CP(clk), .Q(\memory[25][26] ) );
  CFD1QXL \memory_reg[25][25]  ( .D(n572), .CP(clk), .Q(\memory[25][25] ) );
  CFD1QXL \memory_reg[25][24]  ( .D(n573), .CP(clk), .Q(\memory[25][24] ) );
  CFD1QXL \memory_reg[25][23]  ( .D(n574), .CP(clk), .Q(\memory[25][23] ) );
  CFD1QXL \memory_reg[25][22]  ( .D(n575), .CP(clk), .Q(\memory[25][22] ) );
  CFD1QXL \memory_reg[25][21]  ( .D(n576), .CP(clk), .Q(\memory[25][21] ) );
  CFD1QXL \memory_reg[25][20]  ( .D(n577), .CP(clk), .Q(\memory[25][20] ) );
  CFD1QXL \memory_reg[25][19]  ( .D(n578), .CP(clk), .Q(\memory[25][19] ) );
  CFD1QXL \memory_reg[25][18]  ( .D(n579), .CP(clk), .Q(\memory[25][18] ) );
  CFD1QXL \memory_reg[25][17]  ( .D(n580), .CP(clk), .Q(\memory[25][17] ) );
  CFD1QXL \memory_reg[25][16]  ( .D(n581), .CP(clk), .Q(\memory[25][16] ) );
  CFD1QXL \memory_reg[25][15]  ( .D(n582), .CP(clk), .Q(\memory[25][15] ) );
  CFD1QXL \memory_reg[25][14]  ( .D(n583), .CP(clk), .Q(\memory[25][14] ) );
  CFD1QXL \memory_reg[25][13]  ( .D(n584), .CP(clk), .Q(\memory[25][13] ) );
  CFD1QXL \memory_reg[25][12]  ( .D(n585), .CP(clk), .Q(\memory[25][12] ) );
  CFD1QXL \memory_reg[25][11]  ( .D(n586), .CP(clk), .Q(\memory[25][11] ) );
  CFD1QXL \memory_reg[25][10]  ( .D(n587), .CP(clk), .Q(\memory[25][10] ) );
  CFD1QXL \memory_reg[25][9]  ( .D(n588), .CP(clk), .Q(\memory[25][9] ) );
  CFD1QXL \memory_reg[25][8]  ( .D(n589), .CP(clk), .Q(\memory[25][8] ) );
  CFD1QXL \memory_reg[25][7]  ( .D(n590), .CP(clk), .Q(\memory[25][7] ) );
  CFD1QXL \memory_reg[25][6]  ( .D(n591), .CP(clk), .Q(\memory[25][6] ) );
  CFD1QXL \memory_reg[25][5]  ( .D(n592), .CP(clk), .Q(\memory[25][5] ) );
  CFD1QXL \memory_reg[25][4]  ( .D(n593), .CP(clk), .Q(\memory[25][4] ) );
  CFD1QXL \memory_reg[25][3]  ( .D(n594), .CP(clk), .Q(\memory[25][3] ) );
  CFD1QXL \memory_reg[25][2]  ( .D(n595), .CP(clk), .Q(\memory[25][2] ) );
  CFD1QXL \memory_reg[25][1]  ( .D(n596), .CP(clk), .Q(\memory[25][1] ) );
  CFD1QXL \memory_reg[25][0]  ( .D(n597), .CP(clk), .Q(\memory[25][0] ) );
  CFD1QXL \memory_reg[24][63]  ( .D(n605), .CP(clk), .Q(\memory[24][63] ) );
  CFD1QXL \memory_reg[24][62]  ( .D(n606), .CP(clk), .Q(\memory[24][62] ) );
  CFD1QXL \memory_reg[24][61]  ( .D(n607), .CP(clk), .Q(\memory[24][61] ) );
  CFD1QXL \memory_reg[24][60]  ( .D(n608), .CP(clk), .Q(\memory[24][60] ) );
  CFD1QXL \memory_reg[24][59]  ( .D(n609), .CP(clk), .Q(\memory[24][59] ) );
  CFD1QXL \memory_reg[24][58]  ( .D(n610), .CP(clk), .Q(\memory[24][58] ) );
  CFD1QXL \memory_reg[24][57]  ( .D(n611), .CP(clk), .Q(\memory[24][57] ) );
  CFD1QXL \memory_reg[24][56]  ( .D(n612), .CP(clk), .Q(\memory[24][56] ) );
  CFD1QXL \memory_reg[24][55]  ( .D(n613), .CP(clk), .Q(\memory[24][55] ) );
  CFD1QXL \memory_reg[24][54]  ( .D(n614), .CP(clk), .Q(\memory[24][54] ) );
  CFD1QXL \memory_reg[24][53]  ( .D(n615), .CP(clk), .Q(\memory[24][53] ) );
  CFD1QXL \memory_reg[24][52]  ( .D(n616), .CP(clk), .Q(\memory[24][52] ) );
  CFD1QXL \memory_reg[24][51]  ( .D(n617), .CP(clk), .Q(\memory[24][51] ) );
  CFD1QXL \memory_reg[24][50]  ( .D(n618), .CP(clk), .Q(\memory[24][50] ) );
  CFD1QXL \memory_reg[24][49]  ( .D(n619), .CP(clk), .Q(\memory[24][49] ) );
  CFD1QXL \memory_reg[24][48]  ( .D(n620), .CP(clk), .Q(\memory[24][48] ) );
  CFD1QXL \memory_reg[24][47]  ( .D(n621), .CP(clk), .Q(\memory[24][47] ) );
  CFD1QXL \memory_reg[24][46]  ( .D(n622), .CP(clk), .Q(\memory[24][46] ) );
  CFD1QXL \memory_reg[24][45]  ( .D(n623), .CP(clk), .Q(\memory[24][45] ) );
  CFD1QXL \memory_reg[24][44]  ( .D(n624), .CP(clk), .Q(\memory[24][44] ) );
  CFD1QXL \memory_reg[24][43]  ( .D(n625), .CP(clk), .Q(\memory[24][43] ) );
  CFD1QXL \memory_reg[24][42]  ( .D(n626), .CP(clk), .Q(\memory[24][42] ) );
  CFD1QXL \memory_reg[24][41]  ( .D(n627), .CP(clk), .Q(\memory[24][41] ) );
  CFD1QXL \memory_reg[24][40]  ( .D(n628), .CP(clk), .Q(\memory[24][40] ) );
  CFD1QXL \memory_reg[24][39]  ( .D(n629), .CP(clk), .Q(\memory[24][39] ) );
  CFD1QXL \memory_reg[24][38]  ( .D(n630), .CP(clk), .Q(\memory[24][38] ) );
  CFD1QXL \memory_reg[24][37]  ( .D(n631), .CP(clk), .Q(\memory[24][37] ) );
  CFD1QXL \memory_reg[24][36]  ( .D(n632), .CP(clk), .Q(\memory[24][36] ) );
  CFD1QXL \memory_reg[24][35]  ( .D(n633), .CP(clk), .Q(\memory[24][35] ) );
  CFD1QXL \memory_reg[24][34]  ( .D(n634), .CP(clk), .Q(\memory[24][34] ) );
  CFD1QXL \memory_reg[24][33]  ( .D(n635), .CP(clk), .Q(\memory[24][33] ) );
  CFD1QXL \memory_reg[24][32]  ( .D(n636), .CP(clk), .Q(\memory[24][32] ) );
  CFD1QXL \memory_reg[24][31]  ( .D(n637), .CP(clk), .Q(\memory[24][31] ) );
  CFD1QXL \memory_reg[24][30]  ( .D(n638), .CP(clk), .Q(\memory[24][30] ) );
  CFD1QXL \memory_reg[24][29]  ( .D(n639), .CP(clk), .Q(\memory[24][29] ) );
  CFD1QXL \memory_reg[24][28]  ( .D(n640), .CP(clk), .Q(\memory[24][28] ) );
  CFD1QXL \memory_reg[24][27]  ( .D(n641), .CP(clk), .Q(\memory[24][27] ) );
  CFD1QXL \memory_reg[24][26]  ( .D(n642), .CP(clk), .Q(\memory[24][26] ) );
  CFD1QXL \memory_reg[24][25]  ( .D(n643), .CP(clk), .Q(\memory[24][25] ) );
  CFD1QXL \memory_reg[24][24]  ( .D(n644), .CP(clk), .Q(\memory[24][24] ) );
  CFD1QXL \memory_reg[24][23]  ( .D(n645), .CP(clk), .Q(\memory[24][23] ) );
  CFD1QXL \memory_reg[24][22]  ( .D(n646), .CP(clk), .Q(\memory[24][22] ) );
  CFD1QXL \memory_reg[24][21]  ( .D(n647), .CP(clk), .Q(\memory[24][21] ) );
  CFD1QXL \memory_reg[24][20]  ( .D(n648), .CP(clk), .Q(\memory[24][20] ) );
  CFD1QXL \memory_reg[24][19]  ( .D(n649), .CP(clk), .Q(\memory[24][19] ) );
  CFD1QXL \memory_reg[24][18]  ( .D(n650), .CP(clk), .Q(\memory[24][18] ) );
  CFD1QXL \memory_reg[24][17]  ( .D(n651), .CP(clk), .Q(\memory[24][17] ) );
  CFD1QXL \memory_reg[24][16]  ( .D(n652), .CP(clk), .Q(\memory[24][16] ) );
  CFD1QXL \memory_reg[24][15]  ( .D(n653), .CP(clk), .Q(\memory[24][15] ) );
  CFD1QXL \memory_reg[24][14]  ( .D(n654), .CP(clk), .Q(\memory[24][14] ) );
  CFD1QXL \memory_reg[24][13]  ( .D(n655), .CP(clk), .Q(\memory[24][13] ) );
  CFD1QXL \memory_reg[24][12]  ( .D(n656), .CP(clk), .Q(\memory[24][12] ) );
  CFD1QXL \memory_reg[24][11]  ( .D(n657), .CP(clk), .Q(\memory[24][11] ) );
  CFD1QXL \memory_reg[24][10]  ( .D(n658), .CP(clk), .Q(\memory[24][10] ) );
  CFD1QXL \memory_reg[24][9]  ( .D(n659), .CP(clk), .Q(\memory[24][9] ) );
  CFD1QXL \memory_reg[24][8]  ( .D(n660), .CP(clk), .Q(\memory[24][8] ) );
  CFD1QXL \memory_reg[24][7]  ( .D(n661), .CP(clk), .Q(\memory[24][7] ) );
  CFD1QXL \memory_reg[24][6]  ( .D(n662), .CP(clk), .Q(\memory[24][6] ) );
  CFD1QXL \memory_reg[24][5]  ( .D(n663), .CP(clk), .Q(\memory[24][5] ) );
  CFD1QXL \memory_reg[24][4]  ( .D(n664), .CP(clk), .Q(\memory[24][4] ) );
  CFD1QXL \memory_reg[24][3]  ( .D(n665), .CP(clk), .Q(\memory[24][3] ) );
  CFD1QXL \memory_reg[24][2]  ( .D(n666), .CP(clk), .Q(\memory[24][2] ) );
  CFD1QXL \memory_reg[24][1]  ( .D(n667), .CP(clk), .Q(\memory[24][1] ) );
  CFD1QXL \memory_reg[24][0]  ( .D(n668), .CP(clk), .Q(\memory[24][0] ) );
  CFD1QXL \memory_reg[22][63]  ( .D(n747), .CP(clk), .Q(\memory[22][63] ) );
  CFD1QXL \memory_reg[22][62]  ( .D(n748), .CP(clk), .Q(\memory[22][62] ) );
  CFD1QXL \memory_reg[22][61]  ( .D(n749), .CP(clk), .Q(\memory[22][61] ) );
  CFD1QXL \memory_reg[22][60]  ( .D(n750), .CP(clk), .Q(\memory[22][60] ) );
  CFD1QXL \memory_reg[22][59]  ( .D(n751), .CP(clk), .Q(\memory[22][59] ) );
  CFD1QXL \memory_reg[22][58]  ( .D(n752), .CP(clk), .Q(\memory[22][58] ) );
  CFD1QXL \memory_reg[22][57]  ( .D(n753), .CP(clk), .Q(\memory[22][57] ) );
  CFD1QXL \memory_reg[22][56]  ( .D(n754), .CP(clk), .Q(\memory[22][56] ) );
  CFD1QXL \memory_reg[22][55]  ( .D(n755), .CP(clk), .Q(\memory[22][55] ) );
  CFD1QXL \memory_reg[22][54]  ( .D(n756), .CP(clk), .Q(\memory[22][54] ) );
  CFD1QXL \memory_reg[22][53]  ( .D(n757), .CP(clk), .Q(\memory[22][53] ) );
  CFD1QXL \memory_reg[22][52]  ( .D(n758), .CP(clk), .Q(\memory[22][52] ) );
  CFD1QXL \memory_reg[22][51]  ( .D(n759), .CP(clk), .Q(\memory[22][51] ) );
  CFD1QXL \memory_reg[22][50]  ( .D(n760), .CP(clk), .Q(\memory[22][50] ) );
  CFD1QXL \memory_reg[22][49]  ( .D(n761), .CP(clk), .Q(\memory[22][49] ) );
  CFD1QXL \memory_reg[22][48]  ( .D(n762), .CP(clk), .Q(\memory[22][48] ) );
  CFD1QXL \memory_reg[22][47]  ( .D(n763), .CP(clk), .Q(\memory[22][47] ) );
  CFD1QXL \memory_reg[22][46]  ( .D(n764), .CP(clk), .Q(\memory[22][46] ) );
  CFD1QXL \memory_reg[22][45]  ( .D(n765), .CP(clk), .Q(\memory[22][45] ) );
  CFD1QXL \memory_reg[22][44]  ( .D(n766), .CP(clk), .Q(\memory[22][44] ) );
  CFD1QXL \memory_reg[22][43]  ( .D(n767), .CP(clk), .Q(\memory[22][43] ) );
  CFD1QXL \memory_reg[22][42]  ( .D(n768), .CP(clk), .Q(\memory[22][42] ) );
  CFD1QXL \memory_reg[22][41]  ( .D(n769), .CP(clk), .Q(\memory[22][41] ) );
  CFD1QXL \memory_reg[22][40]  ( .D(n770), .CP(clk), .Q(\memory[22][40] ) );
  CFD1QXL \memory_reg[22][39]  ( .D(n771), .CP(clk), .Q(\memory[22][39] ) );
  CFD1QXL \memory_reg[22][38]  ( .D(n772), .CP(clk), .Q(\memory[22][38] ) );
  CFD1QXL \memory_reg[22][37]  ( .D(n773), .CP(clk), .Q(\memory[22][37] ) );
  CFD1QXL \memory_reg[22][36]  ( .D(n774), .CP(clk), .Q(\memory[22][36] ) );
  CFD1QXL \memory_reg[22][35]  ( .D(n775), .CP(clk), .Q(\memory[22][35] ) );
  CFD1QXL \memory_reg[22][34]  ( .D(n776), .CP(clk), .Q(\memory[22][34] ) );
  CFD1QXL \memory_reg[22][33]  ( .D(n777), .CP(clk), .Q(\memory[22][33] ) );
  CFD1QXL \memory_reg[22][32]  ( .D(n778), .CP(clk), .Q(\memory[22][32] ) );
  CFD1QXL \memory_reg[22][31]  ( .D(n779), .CP(clk), .Q(\memory[22][31] ) );
  CFD1QXL \memory_reg[22][30]  ( .D(n780), .CP(clk), .Q(\memory[22][30] ) );
  CFD1QXL \memory_reg[22][29]  ( .D(n781), .CP(clk), .Q(\memory[22][29] ) );
  CFD1QXL \memory_reg[22][28]  ( .D(n782), .CP(clk), .Q(\memory[22][28] ) );
  CFD1QXL \memory_reg[22][27]  ( .D(n783), .CP(clk), .Q(\memory[22][27] ) );
  CFD1QXL \memory_reg[22][26]  ( .D(n784), .CP(clk), .Q(\memory[22][26] ) );
  CFD1QXL \memory_reg[22][25]  ( .D(n785), .CP(clk), .Q(\memory[22][25] ) );
  CFD1QXL \memory_reg[22][24]  ( .D(n786), .CP(clk), .Q(\memory[22][24] ) );
  CFD1QXL \memory_reg[22][23]  ( .D(n787), .CP(clk), .Q(\memory[22][23] ) );
  CFD1QXL \memory_reg[22][22]  ( .D(n788), .CP(clk), .Q(\memory[22][22] ) );
  CFD1QXL \memory_reg[22][21]  ( .D(n789), .CP(clk), .Q(\memory[22][21] ) );
  CFD1QXL \memory_reg[22][20]  ( .D(n790), .CP(clk), .Q(\memory[22][20] ) );
  CFD1QXL \memory_reg[22][19]  ( .D(n791), .CP(clk), .Q(\memory[22][19] ) );
  CFD1QXL \memory_reg[22][18]  ( .D(n792), .CP(clk), .Q(\memory[22][18] ) );
  CFD1QXL \memory_reg[22][17]  ( .D(n793), .CP(clk), .Q(\memory[22][17] ) );
  CFD1QXL \memory_reg[22][16]  ( .D(n794), .CP(clk), .Q(\memory[22][16] ) );
  CFD1QXL \memory_reg[22][15]  ( .D(n795), .CP(clk), .Q(\memory[22][15] ) );
  CFD1QXL \memory_reg[22][14]  ( .D(n796), .CP(clk), .Q(\memory[22][14] ) );
  CFD1QXL \memory_reg[22][13]  ( .D(n797), .CP(clk), .Q(\memory[22][13] ) );
  CFD1QXL \memory_reg[22][12]  ( .D(n798), .CP(clk), .Q(\memory[22][12] ) );
  CFD1QXL \memory_reg[22][11]  ( .D(n799), .CP(clk), .Q(\memory[22][11] ) );
  CFD1QXL \memory_reg[22][10]  ( .D(n800), .CP(clk), .Q(\memory[22][10] ) );
  CFD1QXL \memory_reg[22][9]  ( .D(n801), .CP(clk), .Q(\memory[22][9] ) );
  CFD1QXL \memory_reg[22][8]  ( .D(n802), .CP(clk), .Q(\memory[22][8] ) );
  CFD1QXL \memory_reg[22][7]  ( .D(n803), .CP(clk), .Q(\memory[22][7] ) );
  CFD1QXL \memory_reg[22][6]  ( .D(n804), .CP(clk), .Q(\memory[22][6] ) );
  CFD1QXL \memory_reg[22][5]  ( .D(n805), .CP(clk), .Q(\memory[22][5] ) );
  CFD1QXL \memory_reg[22][4]  ( .D(n806), .CP(clk), .Q(\memory[22][4] ) );
  CFD1QXL \memory_reg[22][3]  ( .D(n807), .CP(clk), .Q(\memory[22][3] ) );
  CFD1QXL \memory_reg[22][2]  ( .D(n808), .CP(clk), .Q(\memory[22][2] ) );
  CFD1QXL \memory_reg[22][1]  ( .D(n809), .CP(clk), .Q(\memory[22][1] ) );
  CFD1QXL \memory_reg[22][0]  ( .D(n810), .CP(clk), .Q(\memory[22][0] ) );
  CFD1QXL \memory_reg[21][63]  ( .D(n818), .CP(clk), .Q(\memory[21][63] ) );
  CFD1QXL \memory_reg[21][62]  ( .D(n819), .CP(clk), .Q(\memory[21][62] ) );
  CFD1QXL \memory_reg[21][61]  ( .D(n820), .CP(clk), .Q(\memory[21][61] ) );
  CFD1QXL \memory_reg[21][60]  ( .D(n821), .CP(clk), .Q(\memory[21][60] ) );
  CFD1QXL \memory_reg[21][59]  ( .D(n822), .CP(clk), .Q(\memory[21][59] ) );
  CFD1QXL \memory_reg[21][58]  ( .D(n823), .CP(clk), .Q(\memory[21][58] ) );
  CFD1QXL \memory_reg[21][57]  ( .D(n824), .CP(clk), .Q(\memory[21][57] ) );
  CFD1QXL \memory_reg[21][56]  ( .D(n825), .CP(clk), .Q(\memory[21][56] ) );
  CFD1QXL \memory_reg[21][55]  ( .D(n826), .CP(clk), .Q(\memory[21][55] ) );
  CFD1QXL \memory_reg[21][54]  ( .D(n827), .CP(clk), .Q(\memory[21][54] ) );
  CFD1QXL \memory_reg[21][53]  ( .D(n828), .CP(clk), .Q(\memory[21][53] ) );
  CFD1QXL \memory_reg[21][52]  ( .D(n829), .CP(clk), .Q(\memory[21][52] ) );
  CFD1QXL \memory_reg[21][51]  ( .D(n830), .CP(clk), .Q(\memory[21][51] ) );
  CFD1QXL \memory_reg[21][50]  ( .D(n831), .CP(clk), .Q(\memory[21][50] ) );
  CFD1QXL \memory_reg[21][49]  ( .D(n832), .CP(clk), .Q(\memory[21][49] ) );
  CFD1QXL \memory_reg[21][48]  ( .D(n833), .CP(clk), .Q(\memory[21][48] ) );
  CFD1QXL \memory_reg[21][47]  ( .D(n834), .CP(clk), .Q(\memory[21][47] ) );
  CFD1QXL \memory_reg[21][46]  ( .D(n835), .CP(clk), .Q(\memory[21][46] ) );
  CFD1QXL \memory_reg[21][45]  ( .D(n836), .CP(clk), .Q(\memory[21][45] ) );
  CFD1QXL \memory_reg[21][44]  ( .D(n837), .CP(clk), .Q(\memory[21][44] ) );
  CFD1QXL \memory_reg[21][43]  ( .D(n838), .CP(clk), .Q(\memory[21][43] ) );
  CFD1QXL \memory_reg[21][42]  ( .D(n839), .CP(clk), .Q(\memory[21][42] ) );
  CFD1QXL \memory_reg[21][41]  ( .D(n840), .CP(clk), .Q(\memory[21][41] ) );
  CFD1QXL \memory_reg[21][40]  ( .D(n841), .CP(clk), .Q(\memory[21][40] ) );
  CFD1QXL \memory_reg[21][39]  ( .D(n842), .CP(clk), .Q(\memory[21][39] ) );
  CFD1QXL \memory_reg[21][38]  ( .D(n843), .CP(clk), .Q(\memory[21][38] ) );
  CFD1QXL \memory_reg[21][37]  ( .D(n844), .CP(clk), .Q(\memory[21][37] ) );
  CFD1QXL \memory_reg[21][36]  ( .D(n845), .CP(clk), .Q(\memory[21][36] ) );
  CFD1QXL \memory_reg[21][35]  ( .D(n846), .CP(clk), .Q(\memory[21][35] ) );
  CFD1QXL \memory_reg[21][34]  ( .D(n847), .CP(clk), .Q(\memory[21][34] ) );
  CFD1QXL \memory_reg[21][33]  ( .D(n848), .CP(clk), .Q(\memory[21][33] ) );
  CFD1QXL \memory_reg[21][32]  ( .D(n849), .CP(clk), .Q(\memory[21][32] ) );
  CFD1QXL \memory_reg[21][31]  ( .D(n850), .CP(clk), .Q(\memory[21][31] ) );
  CFD1QXL \memory_reg[21][30]  ( .D(n851), .CP(clk), .Q(\memory[21][30] ) );
  CFD1QXL \memory_reg[21][29]  ( .D(n852), .CP(clk), .Q(\memory[21][29] ) );
  CFD1QXL \memory_reg[21][28]  ( .D(n853), .CP(clk), .Q(\memory[21][28] ) );
  CFD1QXL \memory_reg[21][27]  ( .D(n854), .CP(clk), .Q(\memory[21][27] ) );
  CFD1QXL \memory_reg[21][26]  ( .D(n855), .CP(clk), .Q(\memory[21][26] ) );
  CFD1QXL \memory_reg[21][25]  ( .D(n856), .CP(clk), .Q(\memory[21][25] ) );
  CFD1QXL \memory_reg[21][24]  ( .D(n857), .CP(clk), .Q(\memory[21][24] ) );
  CFD1QXL \memory_reg[21][23]  ( .D(n858), .CP(clk), .Q(\memory[21][23] ) );
  CFD1QXL \memory_reg[21][22]  ( .D(n859), .CP(clk), .Q(\memory[21][22] ) );
  CFD1QXL \memory_reg[21][21]  ( .D(n860), .CP(clk), .Q(\memory[21][21] ) );
  CFD1QXL \memory_reg[21][20]  ( .D(n861), .CP(clk), .Q(\memory[21][20] ) );
  CFD1QXL \memory_reg[21][19]  ( .D(n862), .CP(clk), .Q(\memory[21][19] ) );
  CFD1QXL \memory_reg[21][18]  ( .D(n863), .CP(clk), .Q(\memory[21][18] ) );
  CFD1QXL \memory_reg[21][17]  ( .D(n864), .CP(clk), .Q(\memory[21][17] ) );
  CFD1QXL \memory_reg[21][16]  ( .D(n865), .CP(clk), .Q(\memory[21][16] ) );
  CFD1QXL \memory_reg[21][15]  ( .D(n866), .CP(clk), .Q(\memory[21][15] ) );
  CFD1QXL \memory_reg[21][14]  ( .D(n867), .CP(clk), .Q(\memory[21][14] ) );
  CFD1QXL \memory_reg[21][13]  ( .D(n868), .CP(clk), .Q(\memory[21][13] ) );
  CFD1QXL \memory_reg[21][12]  ( .D(n869), .CP(clk), .Q(\memory[21][12] ) );
  CFD1QXL \memory_reg[21][11]  ( .D(n870), .CP(clk), .Q(\memory[21][11] ) );
  CFD1QXL \memory_reg[21][10]  ( .D(n871), .CP(clk), .Q(\memory[21][10] ) );
  CFD1QXL \memory_reg[21][9]  ( .D(n872), .CP(clk), .Q(\memory[21][9] ) );
  CFD1QXL \memory_reg[21][8]  ( .D(n873), .CP(clk), .Q(\memory[21][8] ) );
  CFD1QXL \memory_reg[21][7]  ( .D(n874), .CP(clk), .Q(\memory[21][7] ) );
  CFD1QXL \memory_reg[21][6]  ( .D(n875), .CP(clk), .Q(\memory[21][6] ) );
  CFD1QXL \memory_reg[21][5]  ( .D(n876), .CP(clk), .Q(\memory[21][5] ) );
  CFD1QXL \memory_reg[21][4]  ( .D(n877), .CP(clk), .Q(\memory[21][4] ) );
  CFD1QXL \memory_reg[21][3]  ( .D(n878), .CP(clk), .Q(\memory[21][3] ) );
  CFD1QXL \memory_reg[21][2]  ( .D(n879), .CP(clk), .Q(\memory[21][2] ) );
  CFD1QXL \memory_reg[21][1]  ( .D(n880), .CP(clk), .Q(\memory[21][1] ) );
  CFD1QXL \memory_reg[21][0]  ( .D(n881), .CP(clk), .Q(\memory[21][0] ) );
  CFD1QXL \memory_reg[20][63]  ( .D(n889), .CP(clk), .Q(\memory[20][63] ) );
  CFD1QXL \memory_reg[20][62]  ( .D(n890), .CP(clk), .Q(\memory[20][62] ) );
  CFD1QXL \memory_reg[20][61]  ( .D(n891), .CP(clk), .Q(\memory[20][61] ) );
  CFD1QXL \memory_reg[20][60]  ( .D(n892), .CP(clk), .Q(\memory[20][60] ) );
  CFD1QXL \memory_reg[20][59]  ( .D(n893), .CP(clk), .Q(\memory[20][59] ) );
  CFD1QXL \memory_reg[20][58]  ( .D(n894), .CP(clk), .Q(\memory[20][58] ) );
  CFD1QXL \memory_reg[20][57]  ( .D(n895), .CP(clk), .Q(\memory[20][57] ) );
  CFD1QXL \memory_reg[20][56]  ( .D(n896), .CP(clk), .Q(\memory[20][56] ) );
  CFD1QXL \memory_reg[20][55]  ( .D(n897), .CP(clk), .Q(\memory[20][55] ) );
  CFD1QXL \memory_reg[20][54]  ( .D(n898), .CP(clk), .Q(\memory[20][54] ) );
  CFD1QXL \memory_reg[20][53]  ( .D(n899), .CP(clk), .Q(\memory[20][53] ) );
  CFD1QXL \memory_reg[20][52]  ( .D(n900), .CP(clk), .Q(\memory[20][52] ) );
  CFD1QXL \memory_reg[20][51]  ( .D(n901), .CP(clk), .Q(\memory[20][51] ) );
  CFD1QXL \memory_reg[20][50]  ( .D(n902), .CP(clk), .Q(\memory[20][50] ) );
  CFD1QXL \memory_reg[20][49]  ( .D(n903), .CP(clk), .Q(\memory[20][49] ) );
  CFD1QXL \memory_reg[20][48]  ( .D(n904), .CP(clk), .Q(\memory[20][48] ) );
  CFD1QXL \memory_reg[20][47]  ( .D(n905), .CP(clk), .Q(\memory[20][47] ) );
  CFD1QXL \memory_reg[20][46]  ( .D(n906), .CP(clk), .Q(\memory[20][46] ) );
  CFD1QXL \memory_reg[20][45]  ( .D(n907), .CP(clk), .Q(\memory[20][45] ) );
  CFD1QXL \memory_reg[20][44]  ( .D(n908), .CP(clk), .Q(\memory[20][44] ) );
  CFD1QXL \memory_reg[20][43]  ( .D(n909), .CP(clk), .Q(\memory[20][43] ) );
  CFD1QXL \memory_reg[20][42]  ( .D(n910), .CP(clk), .Q(\memory[20][42] ) );
  CFD1QXL \memory_reg[20][41]  ( .D(n911), .CP(clk), .Q(\memory[20][41] ) );
  CFD1QXL \memory_reg[20][40]  ( .D(n912), .CP(clk), .Q(\memory[20][40] ) );
  CFD1QXL \memory_reg[20][39]  ( .D(n913), .CP(clk), .Q(\memory[20][39] ) );
  CFD1QXL \memory_reg[20][38]  ( .D(n914), .CP(clk), .Q(\memory[20][38] ) );
  CFD1QXL \memory_reg[20][37]  ( .D(n915), .CP(clk), .Q(\memory[20][37] ) );
  CFD1QXL \memory_reg[20][36]  ( .D(n916), .CP(clk), .Q(\memory[20][36] ) );
  CFD1QXL \memory_reg[20][35]  ( .D(n917), .CP(clk), .Q(\memory[20][35] ) );
  CFD1QXL \memory_reg[20][34]  ( .D(n918), .CP(clk), .Q(\memory[20][34] ) );
  CFD1QXL \memory_reg[20][33]  ( .D(n919), .CP(clk), .Q(\memory[20][33] ) );
  CFD1QXL \memory_reg[20][32]  ( .D(n920), .CP(clk), .Q(\memory[20][32] ) );
  CFD1QXL \memory_reg[20][31]  ( .D(n921), .CP(clk), .Q(\memory[20][31] ) );
  CFD1QXL \memory_reg[20][30]  ( .D(n922), .CP(clk), .Q(\memory[20][30] ) );
  CFD1QXL \memory_reg[20][29]  ( .D(n923), .CP(clk), .Q(\memory[20][29] ) );
  CFD1QXL \memory_reg[20][28]  ( .D(n924), .CP(clk), .Q(\memory[20][28] ) );
  CFD1QXL \memory_reg[20][27]  ( .D(n925), .CP(clk), .Q(\memory[20][27] ) );
  CFD1QXL \memory_reg[20][26]  ( .D(n926), .CP(clk), .Q(\memory[20][26] ) );
  CFD1QXL \memory_reg[20][25]  ( .D(n927), .CP(clk), .Q(\memory[20][25] ) );
  CFD1QXL \memory_reg[20][24]  ( .D(n928), .CP(clk), .Q(\memory[20][24] ) );
  CFD1QXL \memory_reg[20][23]  ( .D(n929), .CP(clk), .Q(\memory[20][23] ) );
  CFD1QXL \memory_reg[20][22]  ( .D(n930), .CP(clk), .Q(\memory[20][22] ) );
  CFD1QXL \memory_reg[20][21]  ( .D(n931), .CP(clk), .Q(\memory[20][21] ) );
  CFD1QXL \memory_reg[20][20]  ( .D(n932), .CP(clk), .Q(\memory[20][20] ) );
  CFD1QXL \memory_reg[20][19]  ( .D(n933), .CP(clk), .Q(\memory[20][19] ) );
  CFD1QXL \memory_reg[20][18]  ( .D(n934), .CP(clk), .Q(\memory[20][18] ) );
  CFD1QXL \memory_reg[20][17]  ( .D(n935), .CP(clk), .Q(\memory[20][17] ) );
  CFD1QXL \memory_reg[20][16]  ( .D(n936), .CP(clk), .Q(\memory[20][16] ) );
  CFD1QXL \memory_reg[20][15]  ( .D(n937), .CP(clk), .Q(\memory[20][15] ) );
  CFD1QXL \memory_reg[20][14]  ( .D(n938), .CP(clk), .Q(\memory[20][14] ) );
  CFD1QXL \memory_reg[20][13]  ( .D(n939), .CP(clk), .Q(\memory[20][13] ) );
  CFD1QXL \memory_reg[20][12]  ( .D(n940), .CP(clk), .Q(\memory[20][12] ) );
  CFD1QXL \memory_reg[20][11]  ( .D(n941), .CP(clk), .Q(\memory[20][11] ) );
  CFD1QXL \memory_reg[20][10]  ( .D(n942), .CP(clk), .Q(\memory[20][10] ) );
  CFD1QXL \memory_reg[20][9]  ( .D(n943), .CP(clk), .Q(\memory[20][9] ) );
  CFD1QXL \memory_reg[20][8]  ( .D(n944), .CP(clk), .Q(\memory[20][8] ) );
  CFD1QXL \memory_reg[20][7]  ( .D(n945), .CP(clk), .Q(\memory[20][7] ) );
  CFD1QXL \memory_reg[20][6]  ( .D(n946), .CP(clk), .Q(\memory[20][6] ) );
  CFD1QXL \memory_reg[20][5]  ( .D(n947), .CP(clk), .Q(\memory[20][5] ) );
  CFD1QXL \memory_reg[20][4]  ( .D(n948), .CP(clk), .Q(\memory[20][4] ) );
  CFD1QXL \memory_reg[20][3]  ( .D(n949), .CP(clk), .Q(\memory[20][3] ) );
  CFD1QXL \memory_reg[20][2]  ( .D(n950), .CP(clk), .Q(\memory[20][2] ) );
  CFD1QXL \memory_reg[20][1]  ( .D(n951), .CP(clk), .Q(\memory[20][1] ) );
  CFD1QXL \memory_reg[20][0]  ( .D(n952), .CP(clk), .Q(\memory[20][0] ) );
  CFD1QXL \memory_reg[18][63]  ( .D(n1031), .CP(clk), .Q(\memory[18][63] ) );
  CFD1QXL \memory_reg[18][62]  ( .D(n1032), .CP(clk), .Q(\memory[18][62] ) );
  CFD1QXL \memory_reg[18][61]  ( .D(n1033), .CP(clk), .Q(\memory[18][61] ) );
  CFD1QXL \memory_reg[18][60]  ( .D(n1034), .CP(clk), .Q(\memory[18][60] ) );
  CFD1QXL \memory_reg[18][59]  ( .D(n1035), .CP(clk), .Q(\memory[18][59] ) );
  CFD1QXL \memory_reg[18][58]  ( .D(n1036), .CP(clk), .Q(\memory[18][58] ) );
  CFD1QXL \memory_reg[18][57]  ( .D(n1037), .CP(clk), .Q(\memory[18][57] ) );
  CFD1QXL \memory_reg[18][56]  ( .D(n1038), .CP(clk), .Q(\memory[18][56] ) );
  CFD1QXL \memory_reg[18][55]  ( .D(n1039), .CP(clk), .Q(\memory[18][55] ) );
  CFD1QXL \memory_reg[18][54]  ( .D(n1040), .CP(clk), .Q(\memory[18][54] ) );
  CFD1QXL \memory_reg[18][53]  ( .D(n1041), .CP(clk), .Q(\memory[18][53] ) );
  CFD1QXL \memory_reg[18][52]  ( .D(n1042), .CP(clk), .Q(\memory[18][52] ) );
  CFD1QXL \memory_reg[18][51]  ( .D(n1043), .CP(clk), .Q(\memory[18][51] ) );
  CFD1QXL \memory_reg[18][50]  ( .D(n1044), .CP(clk), .Q(\memory[18][50] ) );
  CFD1QXL \memory_reg[18][49]  ( .D(n1045), .CP(clk), .Q(\memory[18][49] ) );
  CFD1QXL \memory_reg[18][48]  ( .D(n1046), .CP(clk), .Q(\memory[18][48] ) );
  CFD1QXL \memory_reg[18][47]  ( .D(n1047), .CP(clk), .Q(\memory[18][47] ) );
  CFD1QXL \memory_reg[18][46]  ( .D(n1048), .CP(clk), .Q(\memory[18][46] ) );
  CFD1QXL \memory_reg[18][45]  ( .D(n1049), .CP(clk), .Q(\memory[18][45] ) );
  CFD1QXL \memory_reg[18][44]  ( .D(n1050), .CP(clk), .Q(\memory[18][44] ) );
  CFD1QXL \memory_reg[18][43]  ( .D(n1051), .CP(clk), .Q(\memory[18][43] ) );
  CFD1QXL \memory_reg[18][42]  ( .D(n1052), .CP(clk), .Q(\memory[18][42] ) );
  CFD1QXL \memory_reg[18][41]  ( .D(n1053), .CP(clk), .Q(\memory[18][41] ) );
  CFD1QXL \memory_reg[18][40]  ( .D(n1054), .CP(clk), .Q(\memory[18][40] ) );
  CFD1QXL \memory_reg[18][39]  ( .D(n1055), .CP(clk), .Q(\memory[18][39] ) );
  CFD1QXL \memory_reg[18][38]  ( .D(n1056), .CP(clk), .Q(\memory[18][38] ) );
  CFD1QXL \memory_reg[18][37]  ( .D(n1057), .CP(clk), .Q(\memory[18][37] ) );
  CFD1QXL \memory_reg[18][36]  ( .D(n1058), .CP(clk), .Q(\memory[18][36] ) );
  CFD1QXL \memory_reg[18][35]  ( .D(n1059), .CP(clk), .Q(\memory[18][35] ) );
  CFD1QXL \memory_reg[18][34]  ( .D(n1060), .CP(clk), .Q(\memory[18][34] ) );
  CFD1QXL \memory_reg[18][33]  ( .D(n1061), .CP(clk), .Q(\memory[18][33] ) );
  CFD1QXL \memory_reg[18][32]  ( .D(n1062), .CP(clk), .Q(\memory[18][32] ) );
  CFD1QXL \memory_reg[18][31]  ( .D(n1063), .CP(clk), .Q(\memory[18][31] ) );
  CFD1QXL \memory_reg[18][30]  ( .D(n1064), .CP(clk), .Q(\memory[18][30] ) );
  CFD1QXL \memory_reg[18][29]  ( .D(n1065), .CP(clk), .Q(\memory[18][29] ) );
  CFD1QXL \memory_reg[18][28]  ( .D(n1066), .CP(clk), .Q(\memory[18][28] ) );
  CFD1QXL \memory_reg[18][27]  ( .D(n1067), .CP(clk), .Q(\memory[18][27] ) );
  CFD1QXL \memory_reg[18][26]  ( .D(n1068), .CP(clk), .Q(\memory[18][26] ) );
  CFD1QXL \memory_reg[18][25]  ( .D(n1069), .CP(clk), .Q(\memory[18][25] ) );
  CFD1QXL \memory_reg[18][24]  ( .D(n1070), .CP(clk), .Q(\memory[18][24] ) );
  CFD1QXL \memory_reg[18][23]  ( .D(n1071), .CP(clk), .Q(\memory[18][23] ) );
  CFD1QXL \memory_reg[18][22]  ( .D(n1072), .CP(clk), .Q(\memory[18][22] ) );
  CFD1QXL \memory_reg[18][21]  ( .D(n1073), .CP(clk), .Q(\memory[18][21] ) );
  CFD1QXL \memory_reg[18][20]  ( .D(n1074), .CP(clk), .Q(\memory[18][20] ) );
  CFD1QXL \memory_reg[18][19]  ( .D(n1075), .CP(clk), .Q(\memory[18][19] ) );
  CFD1QXL \memory_reg[18][18]  ( .D(n1076), .CP(clk), .Q(\memory[18][18] ) );
  CFD1QXL \memory_reg[18][17]  ( .D(n1077), .CP(clk), .Q(\memory[18][17] ) );
  CFD1QXL \memory_reg[18][16]  ( .D(n1078), .CP(clk), .Q(\memory[18][16] ) );
  CFD1QXL \memory_reg[18][15]  ( .D(n1079), .CP(clk), .Q(\memory[18][15] ) );
  CFD1QXL \memory_reg[18][14]  ( .D(n1080), .CP(clk), .Q(\memory[18][14] ) );
  CFD1QXL \memory_reg[18][13]  ( .D(n1081), .CP(clk), .Q(\memory[18][13] ) );
  CFD1QXL \memory_reg[18][12]  ( .D(n1082), .CP(clk), .Q(\memory[18][12] ) );
  CFD1QXL \memory_reg[18][11]  ( .D(n1083), .CP(clk), .Q(\memory[18][11] ) );
  CFD1QXL \memory_reg[18][10]  ( .D(n1084), .CP(clk), .Q(\memory[18][10] ) );
  CFD1QXL \memory_reg[18][9]  ( .D(n1085), .CP(clk), .Q(\memory[18][9] ) );
  CFD1QXL \memory_reg[18][8]  ( .D(n1086), .CP(clk), .Q(\memory[18][8] ) );
  CFD1QXL \memory_reg[18][7]  ( .D(n1087), .CP(clk), .Q(\memory[18][7] ) );
  CFD1QXL \memory_reg[18][6]  ( .D(n1088), .CP(clk), .Q(\memory[18][6] ) );
  CFD1QXL \memory_reg[18][5]  ( .D(n1089), .CP(clk), .Q(\memory[18][5] ) );
  CFD1QXL \memory_reg[18][4]  ( .D(n1090), .CP(clk), .Q(\memory[18][4] ) );
  CFD1QXL \memory_reg[18][3]  ( .D(n1091), .CP(clk), .Q(\memory[18][3] ) );
  CFD1QXL \memory_reg[18][2]  ( .D(n1092), .CP(clk), .Q(\memory[18][2] ) );
  CFD1QXL \memory_reg[18][1]  ( .D(n1093), .CP(clk), .Q(\memory[18][1] ) );
  CFD1QXL \memory_reg[18][0]  ( .D(n1094), .CP(clk), .Q(\memory[18][0] ) );
  CFD1QXL \memory_reg[17][63]  ( .D(n1102), .CP(clk), .Q(\memory[17][63] ) );
  CFD1QXL \memory_reg[17][62]  ( .D(n1103), .CP(clk), .Q(\memory[17][62] ) );
  CFD1QXL \memory_reg[17][61]  ( .D(n1104), .CP(clk), .Q(\memory[17][61] ) );
  CFD1QXL \memory_reg[17][60]  ( .D(n1105), .CP(clk), .Q(\memory[17][60] ) );
  CFD1QXL \memory_reg[17][59]  ( .D(n1106), .CP(clk), .Q(\memory[17][59] ) );
  CFD1QXL \memory_reg[17][58]  ( .D(n1107), .CP(clk), .Q(\memory[17][58] ) );
  CFD1QXL \memory_reg[17][57]  ( .D(n1108), .CP(clk), .Q(\memory[17][57] ) );
  CFD1QXL \memory_reg[17][56]  ( .D(n1109), .CP(clk), .Q(\memory[17][56] ) );
  CFD1QXL \memory_reg[17][55]  ( .D(n1110), .CP(clk), .Q(\memory[17][55] ) );
  CFD1QXL \memory_reg[17][54]  ( .D(n1111), .CP(clk), .Q(\memory[17][54] ) );
  CFD1QXL \memory_reg[17][53]  ( .D(n1112), .CP(clk), .Q(\memory[17][53] ) );
  CFD1QXL \memory_reg[17][52]  ( .D(n1113), .CP(clk), .Q(\memory[17][52] ) );
  CFD1QXL \memory_reg[17][51]  ( .D(n1114), .CP(clk), .Q(\memory[17][51] ) );
  CFD1QXL \memory_reg[17][50]  ( .D(n1115), .CP(clk), .Q(\memory[17][50] ) );
  CFD1QXL \memory_reg[17][49]  ( .D(n1116), .CP(clk), .Q(\memory[17][49] ) );
  CFD1QXL \memory_reg[17][48]  ( .D(n1117), .CP(clk), .Q(\memory[17][48] ) );
  CFD1QXL \memory_reg[17][47]  ( .D(n1118), .CP(clk), .Q(\memory[17][47] ) );
  CFD1QXL \memory_reg[17][46]  ( .D(n1119), .CP(clk), .Q(\memory[17][46] ) );
  CFD1QXL \memory_reg[17][45]  ( .D(n1120), .CP(clk), .Q(\memory[17][45] ) );
  CFD1QXL \memory_reg[17][44]  ( .D(n1121), .CP(clk), .Q(\memory[17][44] ) );
  CFD1QXL \memory_reg[17][43]  ( .D(n1122), .CP(clk), .Q(\memory[17][43] ) );
  CFD1QXL \memory_reg[17][42]  ( .D(n1123), .CP(clk), .Q(\memory[17][42] ) );
  CFD1QXL \memory_reg[17][41]  ( .D(n1124), .CP(clk), .Q(\memory[17][41] ) );
  CFD1QXL \memory_reg[17][40]  ( .D(n1125), .CP(clk), .Q(\memory[17][40] ) );
  CFD1QXL \memory_reg[17][39]  ( .D(n1126), .CP(clk), .Q(\memory[17][39] ) );
  CFD1QXL \memory_reg[17][38]  ( .D(n1127), .CP(clk), .Q(\memory[17][38] ) );
  CFD1QXL \memory_reg[17][37]  ( .D(n1128), .CP(clk), .Q(\memory[17][37] ) );
  CFD1QXL \memory_reg[17][36]  ( .D(n1129), .CP(clk), .Q(\memory[17][36] ) );
  CFD1QXL \memory_reg[17][35]  ( .D(n1130), .CP(clk), .Q(\memory[17][35] ) );
  CFD1QXL \memory_reg[17][34]  ( .D(n1131), .CP(clk), .Q(\memory[17][34] ) );
  CFD1QXL \memory_reg[17][33]  ( .D(n1132), .CP(clk), .Q(\memory[17][33] ) );
  CFD1QXL \memory_reg[17][32]  ( .D(n1133), .CP(clk), .Q(\memory[17][32] ) );
  CFD1QXL \memory_reg[17][31]  ( .D(n1134), .CP(clk), .Q(\memory[17][31] ) );
  CFD1QXL \memory_reg[17][30]  ( .D(n1135), .CP(clk), .Q(\memory[17][30] ) );
  CFD1QXL \memory_reg[17][29]  ( .D(n1136), .CP(clk), .Q(\memory[17][29] ) );
  CFD1QXL \memory_reg[17][28]  ( .D(n1137), .CP(clk), .Q(\memory[17][28] ) );
  CFD1QXL \memory_reg[17][27]  ( .D(n1138), .CP(clk), .Q(\memory[17][27] ) );
  CFD1QXL \memory_reg[17][26]  ( .D(n1139), .CP(clk), .Q(\memory[17][26] ) );
  CFD1QXL \memory_reg[17][25]  ( .D(n1140), .CP(clk), .Q(\memory[17][25] ) );
  CFD1QXL \memory_reg[17][24]  ( .D(n1141), .CP(clk), .Q(\memory[17][24] ) );
  CFD1QXL \memory_reg[17][23]  ( .D(n1142), .CP(clk), .Q(\memory[17][23] ) );
  CFD1QXL \memory_reg[17][22]  ( .D(n1143), .CP(clk), .Q(\memory[17][22] ) );
  CFD1QXL \memory_reg[17][21]  ( .D(n1144), .CP(clk), .Q(\memory[17][21] ) );
  CFD1QXL \memory_reg[17][20]  ( .D(n1145), .CP(clk), .Q(\memory[17][20] ) );
  CFD1QXL \memory_reg[17][19]  ( .D(n1146), .CP(clk), .Q(\memory[17][19] ) );
  CFD1QXL \memory_reg[17][18]  ( .D(n1147), .CP(clk), .Q(\memory[17][18] ) );
  CFD1QXL \memory_reg[17][17]  ( .D(n1148), .CP(clk), .Q(\memory[17][17] ) );
  CFD1QXL \memory_reg[17][16]  ( .D(n1149), .CP(clk), .Q(\memory[17][16] ) );
  CFD1QXL \memory_reg[17][15]  ( .D(n1150), .CP(clk), .Q(\memory[17][15] ) );
  CFD1QXL \memory_reg[17][14]  ( .D(n1151), .CP(clk), .Q(\memory[17][14] ) );
  CFD1QXL \memory_reg[17][13]  ( .D(n1152), .CP(clk), .Q(\memory[17][13] ) );
  CFD1QXL \memory_reg[17][12]  ( .D(n1153), .CP(clk), .Q(\memory[17][12] ) );
  CFD1QXL \memory_reg[17][11]  ( .D(n1154), .CP(clk), .Q(\memory[17][11] ) );
  CFD1QXL \memory_reg[17][10]  ( .D(n1155), .CP(clk), .Q(\memory[17][10] ) );
  CFD1QXL \memory_reg[17][9]  ( .D(n1156), .CP(clk), .Q(\memory[17][9] ) );
  CFD1QXL \memory_reg[17][8]  ( .D(n1157), .CP(clk), .Q(\memory[17][8] ) );
  CFD1QXL \memory_reg[17][7]  ( .D(n1158), .CP(clk), .Q(\memory[17][7] ) );
  CFD1QXL \memory_reg[17][6]  ( .D(n1159), .CP(clk), .Q(\memory[17][6] ) );
  CFD1QXL \memory_reg[17][5]  ( .D(n1160), .CP(clk), .Q(\memory[17][5] ) );
  CFD1QXL \memory_reg[17][4]  ( .D(n1161), .CP(clk), .Q(\memory[17][4] ) );
  CFD1QXL \memory_reg[17][3]  ( .D(n1162), .CP(clk), .Q(\memory[17][3] ) );
  CFD1QXL \memory_reg[17][2]  ( .D(n1163), .CP(clk), .Q(\memory[17][2] ) );
  CFD1QXL \memory_reg[17][1]  ( .D(n1164), .CP(clk), .Q(\memory[17][1] ) );
  CFD1QXL \memory_reg[17][0]  ( .D(n1165), .CP(clk), .Q(\memory[17][0] ) );
  CFD1QXL \memory_reg[16][63]  ( .D(n1173), .CP(clk), .Q(\memory[16][63] ) );
  CFD1QXL \memory_reg[16][62]  ( .D(n1174), .CP(clk), .Q(\memory[16][62] ) );
  CFD1QXL \memory_reg[16][61]  ( .D(n1175), .CP(clk), .Q(\memory[16][61] ) );
  CFD1QXL \memory_reg[16][60]  ( .D(n1176), .CP(clk), .Q(\memory[16][60] ) );
  CFD1QXL \memory_reg[16][59]  ( .D(n1177), .CP(clk), .Q(\memory[16][59] ) );
  CFD1QXL \memory_reg[16][58]  ( .D(n1178), .CP(clk), .Q(\memory[16][58] ) );
  CFD1QXL \memory_reg[16][57]  ( .D(n1179), .CP(clk), .Q(\memory[16][57] ) );
  CFD1QXL \memory_reg[16][56]  ( .D(n1180), .CP(clk), .Q(\memory[16][56] ) );
  CFD1QXL \memory_reg[16][55]  ( .D(n1181), .CP(clk), .Q(\memory[16][55] ) );
  CFD1QXL \memory_reg[16][54]  ( .D(n1182), .CP(clk), .Q(\memory[16][54] ) );
  CFD1QXL \memory_reg[16][53]  ( .D(n1183), .CP(clk), .Q(\memory[16][53] ) );
  CFD1QXL \memory_reg[16][52]  ( .D(n1184), .CP(clk), .Q(\memory[16][52] ) );
  CFD1QXL \memory_reg[16][51]  ( .D(n1185), .CP(clk), .Q(\memory[16][51] ) );
  CFD1QXL \memory_reg[16][50]  ( .D(n1186), .CP(clk), .Q(\memory[16][50] ) );
  CFD1QXL \memory_reg[16][49]  ( .D(n1187), .CP(clk), .Q(\memory[16][49] ) );
  CFD1QXL \memory_reg[16][48]  ( .D(n1188), .CP(clk), .Q(\memory[16][48] ) );
  CFD1QXL \memory_reg[16][47]  ( .D(n1189), .CP(clk), .Q(\memory[16][47] ) );
  CFD1QXL \memory_reg[16][46]  ( .D(n1190), .CP(clk), .Q(\memory[16][46] ) );
  CFD1QXL \memory_reg[16][45]  ( .D(n1191), .CP(clk), .Q(\memory[16][45] ) );
  CFD1QXL \memory_reg[16][44]  ( .D(n1192), .CP(clk), .Q(\memory[16][44] ) );
  CFD1QXL \memory_reg[16][43]  ( .D(n1193), .CP(clk), .Q(\memory[16][43] ) );
  CFD1QXL \memory_reg[16][42]  ( .D(n1194), .CP(clk), .Q(\memory[16][42] ) );
  CFD1QXL \memory_reg[16][41]  ( .D(n1195), .CP(clk), .Q(\memory[16][41] ) );
  CFD1QXL \memory_reg[16][40]  ( .D(n1196), .CP(clk), .Q(\memory[16][40] ) );
  CFD1QXL \memory_reg[16][39]  ( .D(n1197), .CP(clk), .Q(\memory[16][39] ) );
  CFD1QXL \memory_reg[16][38]  ( .D(n1198), .CP(clk), .Q(\memory[16][38] ) );
  CFD1QXL \memory_reg[16][37]  ( .D(n1199), .CP(clk), .Q(\memory[16][37] ) );
  CFD1QXL \memory_reg[16][36]  ( .D(n1200), .CP(clk), .Q(\memory[16][36] ) );
  CFD1QXL \memory_reg[16][35]  ( .D(n1201), .CP(clk), .Q(\memory[16][35] ) );
  CFD1QXL \memory_reg[16][34]  ( .D(n1202), .CP(clk), .Q(\memory[16][34] ) );
  CFD1QXL \memory_reg[16][33]  ( .D(n1203), .CP(clk), .Q(\memory[16][33] ) );
  CFD1QXL \memory_reg[16][32]  ( .D(n1204), .CP(clk), .Q(\memory[16][32] ) );
  CFD1QXL \memory_reg[16][31]  ( .D(n1205), .CP(clk), .Q(\memory[16][31] ) );
  CFD1QXL \memory_reg[16][30]  ( .D(n1206), .CP(clk), .Q(\memory[16][30] ) );
  CFD1QXL \memory_reg[16][29]  ( .D(n1207), .CP(clk), .Q(\memory[16][29] ) );
  CFD1QXL \memory_reg[16][28]  ( .D(n1208), .CP(clk), .Q(\memory[16][28] ) );
  CFD1QXL \memory_reg[16][27]  ( .D(n1209), .CP(clk), .Q(\memory[16][27] ) );
  CFD1QXL \memory_reg[16][26]  ( .D(n1210), .CP(clk), .Q(\memory[16][26] ) );
  CFD1QXL \memory_reg[16][25]  ( .D(n1211), .CP(clk), .Q(\memory[16][25] ) );
  CFD1QXL \memory_reg[16][24]  ( .D(n1212), .CP(clk), .Q(\memory[16][24] ) );
  CFD1QXL \memory_reg[16][23]  ( .D(n1213), .CP(clk), .Q(\memory[16][23] ) );
  CFD1QXL \memory_reg[16][22]  ( .D(n1214), .CP(clk), .Q(\memory[16][22] ) );
  CFD1QXL \memory_reg[16][21]  ( .D(n1215), .CP(clk), .Q(\memory[16][21] ) );
  CFD1QXL \memory_reg[16][20]  ( .D(n1216), .CP(clk), .Q(\memory[16][20] ) );
  CFD1QXL \memory_reg[16][19]  ( .D(n1217), .CP(clk), .Q(\memory[16][19] ) );
  CFD1QXL \memory_reg[16][18]  ( .D(n1218), .CP(clk), .Q(\memory[16][18] ) );
  CFD1QXL \memory_reg[16][17]  ( .D(n1219), .CP(clk), .Q(\memory[16][17] ) );
  CFD1QXL \memory_reg[16][16]  ( .D(n1220), .CP(clk), .Q(\memory[16][16] ) );
  CFD1QXL \memory_reg[16][15]  ( .D(n1221), .CP(clk), .Q(\memory[16][15] ) );
  CFD1QXL \memory_reg[16][14]  ( .D(n1222), .CP(clk), .Q(\memory[16][14] ) );
  CFD1QXL \memory_reg[16][13]  ( .D(n1223), .CP(clk), .Q(\memory[16][13] ) );
  CFD1QXL \memory_reg[16][12]  ( .D(n1224), .CP(clk), .Q(\memory[16][12] ) );
  CFD1QXL \memory_reg[16][11]  ( .D(n1225), .CP(clk), .Q(\memory[16][11] ) );
  CFD1QXL \memory_reg[16][10]  ( .D(n1226), .CP(clk), .Q(\memory[16][10] ) );
  CFD1QXL \memory_reg[16][9]  ( .D(n1227), .CP(clk), .Q(\memory[16][9] ) );
  CFD1QXL \memory_reg[16][8]  ( .D(n1228), .CP(clk), .Q(\memory[16][8] ) );
  CFD1QXL \memory_reg[16][7]  ( .D(n1229), .CP(clk), .Q(\memory[16][7] ) );
  CFD1QXL \memory_reg[16][6]  ( .D(n1230), .CP(clk), .Q(\memory[16][6] ) );
  CFD1QXL \memory_reg[16][5]  ( .D(n1231), .CP(clk), .Q(\memory[16][5] ) );
  CFD1QXL \memory_reg[16][4]  ( .D(n1232), .CP(clk), .Q(\memory[16][4] ) );
  CFD1QXL \memory_reg[16][3]  ( .D(n1233), .CP(clk), .Q(\memory[16][3] ) );
  CFD1QXL \memory_reg[16][2]  ( .D(n1234), .CP(clk), .Q(\memory[16][2] ) );
  CFD1QXL \memory_reg[16][1]  ( .D(n1235), .CP(clk), .Q(\memory[16][1] ) );
  CFD1QXL \memory_reg[16][0]  ( .D(n1236), .CP(clk), .Q(\memory[16][0] ) );
  CFD1QXL \memory_reg[14][63]  ( .D(n1315), .CP(clk), .Q(\memory[14][63] ) );
  CFD1QXL \memory_reg[14][62]  ( .D(n1316), .CP(clk), .Q(\memory[14][62] ) );
  CFD1QXL \memory_reg[14][61]  ( .D(n1317), .CP(clk), .Q(\memory[14][61] ) );
  CFD1QXL \memory_reg[14][60]  ( .D(n1318), .CP(clk), .Q(\memory[14][60] ) );
  CFD1QXL \memory_reg[14][59]  ( .D(n1319), .CP(clk), .Q(\memory[14][59] ) );
  CFD1QXL \memory_reg[14][58]  ( .D(n1320), .CP(clk), .Q(\memory[14][58] ) );
  CFD1QXL \memory_reg[14][57]  ( .D(n1321), .CP(clk), .Q(\memory[14][57] ) );
  CFD1QXL \memory_reg[14][56]  ( .D(n1322), .CP(clk), .Q(\memory[14][56] ) );
  CFD1QXL \memory_reg[14][55]  ( .D(n1323), .CP(clk), .Q(\memory[14][55] ) );
  CFD1QXL \memory_reg[14][54]  ( .D(n1324), .CP(clk), .Q(\memory[14][54] ) );
  CFD1QXL \memory_reg[14][53]  ( .D(n1325), .CP(clk), .Q(\memory[14][53] ) );
  CFD1QXL \memory_reg[14][52]  ( .D(n1326), .CP(clk), .Q(\memory[14][52] ) );
  CFD1QXL \memory_reg[14][51]  ( .D(n1327), .CP(clk), .Q(\memory[14][51] ) );
  CFD1QXL \memory_reg[14][50]  ( .D(n1328), .CP(clk), .Q(\memory[14][50] ) );
  CFD1QXL \memory_reg[14][49]  ( .D(n1329), .CP(clk), .Q(\memory[14][49] ) );
  CFD1QXL \memory_reg[14][48]  ( .D(n1330), .CP(clk), .Q(\memory[14][48] ) );
  CFD1QXL \memory_reg[14][47]  ( .D(n1331), .CP(clk), .Q(\memory[14][47] ) );
  CFD1QXL \memory_reg[14][46]  ( .D(n1332), .CP(clk), .Q(\memory[14][46] ) );
  CFD1QXL \memory_reg[14][45]  ( .D(n1333), .CP(clk), .Q(\memory[14][45] ) );
  CFD1QXL \memory_reg[14][44]  ( .D(n1334), .CP(clk), .Q(\memory[14][44] ) );
  CFD1QXL \memory_reg[14][43]  ( .D(n1335), .CP(clk), .Q(\memory[14][43] ) );
  CFD1QXL \memory_reg[14][42]  ( .D(n1336), .CP(clk), .Q(\memory[14][42] ) );
  CFD1QXL \memory_reg[14][41]  ( .D(n1337), .CP(clk), .Q(\memory[14][41] ) );
  CFD1QXL \memory_reg[14][40]  ( .D(n1338), .CP(clk), .Q(\memory[14][40] ) );
  CFD1QXL \memory_reg[14][39]  ( .D(n1339), .CP(clk), .Q(\memory[14][39] ) );
  CFD1QXL \memory_reg[14][38]  ( .D(n1340), .CP(clk), .Q(\memory[14][38] ) );
  CFD1QXL \memory_reg[14][37]  ( .D(n1341), .CP(clk), .Q(\memory[14][37] ) );
  CFD1QXL \memory_reg[14][36]  ( .D(n1342), .CP(clk), .Q(\memory[14][36] ) );
  CFD1QXL \memory_reg[14][35]  ( .D(n1343), .CP(clk), .Q(\memory[14][35] ) );
  CFD1QXL \memory_reg[14][34]  ( .D(n1344), .CP(clk), .Q(\memory[14][34] ) );
  CFD1QXL \memory_reg[14][33]  ( .D(n1345), .CP(clk), .Q(\memory[14][33] ) );
  CFD1QXL \memory_reg[14][32]  ( .D(n1346), .CP(clk), .Q(\memory[14][32] ) );
  CFD1QXL \memory_reg[14][31]  ( .D(n1347), .CP(clk), .Q(\memory[14][31] ) );
  CFD1QXL \memory_reg[14][30]  ( .D(n1348), .CP(clk), .Q(\memory[14][30] ) );
  CFD1QXL \memory_reg[14][29]  ( .D(n1349), .CP(clk), .Q(\memory[14][29] ) );
  CFD1QXL \memory_reg[14][28]  ( .D(n1350), .CP(clk), .Q(\memory[14][28] ) );
  CFD1QXL \memory_reg[14][27]  ( .D(n1351), .CP(clk), .Q(\memory[14][27] ) );
  CFD1QXL \memory_reg[14][26]  ( .D(n1352), .CP(clk), .Q(\memory[14][26] ) );
  CFD1QXL \memory_reg[14][25]  ( .D(n1353), .CP(clk), .Q(\memory[14][25] ) );
  CFD1QXL \memory_reg[14][24]  ( .D(n1354), .CP(clk), .Q(\memory[14][24] ) );
  CFD1QXL \memory_reg[14][23]  ( .D(n1355), .CP(clk), .Q(\memory[14][23] ) );
  CFD1QXL \memory_reg[14][22]  ( .D(n1356), .CP(clk), .Q(\memory[14][22] ) );
  CFD1QXL \memory_reg[14][21]  ( .D(n1357), .CP(clk), .Q(\memory[14][21] ) );
  CFD1QXL \memory_reg[14][20]  ( .D(n1358), .CP(clk), .Q(\memory[14][20] ) );
  CFD1QXL \memory_reg[14][19]  ( .D(n1359), .CP(clk), .Q(\memory[14][19] ) );
  CFD1QXL \memory_reg[14][18]  ( .D(n1360), .CP(clk), .Q(\memory[14][18] ) );
  CFD1QXL \memory_reg[14][17]  ( .D(n1361), .CP(clk), .Q(\memory[14][17] ) );
  CFD1QXL \memory_reg[14][16]  ( .D(n1362), .CP(clk), .Q(\memory[14][16] ) );
  CFD1QXL \memory_reg[14][15]  ( .D(n1363), .CP(clk), .Q(\memory[14][15] ) );
  CFD1QXL \memory_reg[14][14]  ( .D(n1364), .CP(clk), .Q(\memory[14][14] ) );
  CFD1QXL \memory_reg[14][13]  ( .D(n1365), .CP(clk), .Q(\memory[14][13] ) );
  CFD1QXL \memory_reg[14][12]  ( .D(n1366), .CP(clk), .Q(\memory[14][12] ) );
  CFD1QXL \memory_reg[14][11]  ( .D(n1367), .CP(clk), .Q(\memory[14][11] ) );
  CFD1QXL \memory_reg[14][10]  ( .D(n1368), .CP(clk), .Q(\memory[14][10] ) );
  CFD1QXL \memory_reg[14][9]  ( .D(n1369), .CP(clk), .Q(\memory[14][9] ) );
  CFD1QXL \memory_reg[14][8]  ( .D(n1370), .CP(clk), .Q(\memory[14][8] ) );
  CFD1QXL \memory_reg[14][7]  ( .D(n1371), .CP(clk), .Q(\memory[14][7] ) );
  CFD1QXL \memory_reg[14][6]  ( .D(n1372), .CP(clk), .Q(\memory[14][6] ) );
  CFD1QXL \memory_reg[14][5]  ( .D(n1373), .CP(clk), .Q(\memory[14][5] ) );
  CFD1QXL \memory_reg[14][4]  ( .D(n1374), .CP(clk), .Q(\memory[14][4] ) );
  CFD1QXL \memory_reg[14][3]  ( .D(n1375), .CP(clk), .Q(\memory[14][3] ) );
  CFD1QXL \memory_reg[14][2]  ( .D(n1376), .CP(clk), .Q(\memory[14][2] ) );
  CFD1QXL \memory_reg[14][1]  ( .D(n1377), .CP(clk), .Q(\memory[14][1] ) );
  CFD1QXL \memory_reg[14][0]  ( .D(n1378), .CP(clk), .Q(\memory[14][0] ) );
  CFD1QXL \memory_reg[13][63]  ( .D(n1386), .CP(clk), .Q(\memory[13][63] ) );
  CFD1QXL \memory_reg[13][62]  ( .D(n1387), .CP(clk), .Q(\memory[13][62] ) );
  CFD1QXL \memory_reg[13][61]  ( .D(n1388), .CP(clk), .Q(\memory[13][61] ) );
  CFD1QXL \memory_reg[13][60]  ( .D(n1389), .CP(clk), .Q(\memory[13][60] ) );
  CFD1QXL \memory_reg[13][59]  ( .D(n1390), .CP(clk), .Q(\memory[13][59] ) );
  CFD1QXL \memory_reg[13][58]  ( .D(n1391), .CP(clk), .Q(\memory[13][58] ) );
  CFD1QXL \memory_reg[13][57]  ( .D(n1392), .CP(clk), .Q(\memory[13][57] ) );
  CFD1QXL \memory_reg[13][56]  ( .D(n1393), .CP(clk), .Q(\memory[13][56] ) );
  CFD1QXL \memory_reg[13][55]  ( .D(n1394), .CP(clk), .Q(\memory[13][55] ) );
  CFD1QXL \memory_reg[13][54]  ( .D(n1395), .CP(clk), .Q(\memory[13][54] ) );
  CFD1QXL \memory_reg[13][53]  ( .D(n1396), .CP(clk), .Q(\memory[13][53] ) );
  CFD1QXL \memory_reg[13][52]  ( .D(n1397), .CP(clk), .Q(\memory[13][52] ) );
  CFD1QXL \memory_reg[13][51]  ( .D(n1398), .CP(clk), .Q(\memory[13][51] ) );
  CFD1QXL \memory_reg[13][50]  ( .D(n1399), .CP(clk), .Q(\memory[13][50] ) );
  CFD1QXL \memory_reg[13][49]  ( .D(n1400), .CP(clk), .Q(\memory[13][49] ) );
  CFD1QXL \memory_reg[13][48]  ( .D(n1401), .CP(clk), .Q(\memory[13][48] ) );
  CFD1QXL \memory_reg[13][47]  ( .D(n1402), .CP(clk), .Q(\memory[13][47] ) );
  CFD1QXL \memory_reg[13][46]  ( .D(n1403), .CP(clk), .Q(\memory[13][46] ) );
  CFD1QXL \memory_reg[13][45]  ( .D(n1404), .CP(clk), .Q(\memory[13][45] ) );
  CFD1QXL \memory_reg[13][44]  ( .D(n1405), .CP(clk), .Q(\memory[13][44] ) );
  CFD1QXL \memory_reg[13][43]  ( .D(n1406), .CP(clk), .Q(\memory[13][43] ) );
  CFD1QXL \memory_reg[13][42]  ( .D(n1407), .CP(clk), .Q(\memory[13][42] ) );
  CFD1QXL \memory_reg[13][41]  ( .D(n1408), .CP(clk), .Q(\memory[13][41] ) );
  CFD1QXL \memory_reg[13][40]  ( .D(n1409), .CP(clk), .Q(\memory[13][40] ) );
  CFD1QXL \memory_reg[13][39]  ( .D(n1410), .CP(clk), .Q(\memory[13][39] ) );
  CFD1QXL \memory_reg[13][38]  ( .D(n1411), .CP(clk), .Q(\memory[13][38] ) );
  CFD1QXL \memory_reg[13][37]  ( .D(n1412), .CP(clk), .Q(\memory[13][37] ) );
  CFD1QXL \memory_reg[13][36]  ( .D(n1413), .CP(clk), .Q(\memory[13][36] ) );
  CFD1QXL \memory_reg[13][35]  ( .D(n1414), .CP(clk), .Q(\memory[13][35] ) );
  CFD1QXL \memory_reg[13][34]  ( .D(n1415), .CP(clk), .Q(\memory[13][34] ) );
  CFD1QXL \memory_reg[13][33]  ( .D(n1416), .CP(clk), .Q(\memory[13][33] ) );
  CFD1QXL \memory_reg[13][32]  ( .D(n1417), .CP(clk), .Q(\memory[13][32] ) );
  CFD1QXL \memory_reg[13][31]  ( .D(n1418), .CP(clk), .Q(\memory[13][31] ) );
  CFD1QXL \memory_reg[13][30]  ( .D(n1419), .CP(clk), .Q(\memory[13][30] ) );
  CFD1QXL \memory_reg[13][29]  ( .D(n1420), .CP(clk), .Q(\memory[13][29] ) );
  CFD1QXL \memory_reg[13][28]  ( .D(n1421), .CP(clk), .Q(\memory[13][28] ) );
  CFD1QXL \memory_reg[13][27]  ( .D(n1422), .CP(clk), .Q(\memory[13][27] ) );
  CFD1QXL \memory_reg[13][26]  ( .D(n1423), .CP(clk), .Q(\memory[13][26] ) );
  CFD1QXL \memory_reg[13][25]  ( .D(n1424), .CP(clk), .Q(\memory[13][25] ) );
  CFD1QXL \memory_reg[13][24]  ( .D(n1425), .CP(clk), .Q(\memory[13][24] ) );
  CFD1QXL \memory_reg[13][23]  ( .D(n1426), .CP(clk), .Q(\memory[13][23] ) );
  CFD1QXL \memory_reg[13][22]  ( .D(n1427), .CP(clk), .Q(\memory[13][22] ) );
  CFD1QXL \memory_reg[13][21]  ( .D(n1428), .CP(clk), .Q(\memory[13][21] ) );
  CFD1QXL \memory_reg[13][20]  ( .D(n1429), .CP(clk), .Q(\memory[13][20] ) );
  CFD1QXL \memory_reg[13][19]  ( .D(n1430), .CP(clk), .Q(\memory[13][19] ) );
  CFD1QXL \memory_reg[13][18]  ( .D(n1431), .CP(clk), .Q(\memory[13][18] ) );
  CFD1QXL \memory_reg[13][17]  ( .D(n1432), .CP(clk), .Q(\memory[13][17] ) );
  CFD1QXL \memory_reg[13][16]  ( .D(n1433), .CP(clk), .Q(\memory[13][16] ) );
  CFD1QXL \memory_reg[13][15]  ( .D(n1434), .CP(clk), .Q(\memory[13][15] ) );
  CFD1QXL \memory_reg[13][14]  ( .D(n1435), .CP(clk), .Q(\memory[13][14] ) );
  CFD1QXL \memory_reg[13][13]  ( .D(n1436), .CP(clk), .Q(\memory[13][13] ) );
  CFD1QXL \memory_reg[13][12]  ( .D(n1437), .CP(clk), .Q(\memory[13][12] ) );
  CFD1QXL \memory_reg[13][11]  ( .D(n1438), .CP(clk), .Q(\memory[13][11] ) );
  CFD1QXL \memory_reg[13][10]  ( .D(n1439), .CP(clk), .Q(\memory[13][10] ) );
  CFD1QXL \memory_reg[13][9]  ( .D(n1440), .CP(clk), .Q(\memory[13][9] ) );
  CFD1QXL \memory_reg[13][8]  ( .D(n1441), .CP(clk), .Q(\memory[13][8] ) );
  CFD1QXL \memory_reg[13][7]  ( .D(n1442), .CP(clk), .Q(\memory[13][7] ) );
  CFD1QXL \memory_reg[13][6]  ( .D(n1443), .CP(clk), .Q(\memory[13][6] ) );
  CFD1QXL \memory_reg[13][5]  ( .D(n1444), .CP(clk), .Q(\memory[13][5] ) );
  CFD1QXL \memory_reg[13][4]  ( .D(n1445), .CP(clk), .Q(\memory[13][4] ) );
  CFD1QXL \memory_reg[13][3]  ( .D(n1446), .CP(clk), .Q(\memory[13][3] ) );
  CFD1QXL \memory_reg[13][2]  ( .D(n1447), .CP(clk), .Q(\memory[13][2] ) );
  CFD1QXL \memory_reg[13][1]  ( .D(n1448), .CP(clk), .Q(\memory[13][1] ) );
  CFD1QXL \memory_reg[13][0]  ( .D(n1449), .CP(clk), .Q(\memory[13][0] ) );
  CFD1QXL \memory_reg[12][63]  ( .D(n1457), .CP(clk), .Q(\memory[12][63] ) );
  CFD1QXL \memory_reg[12][62]  ( .D(n1458), .CP(clk), .Q(\memory[12][62] ) );
  CFD1QXL \memory_reg[12][61]  ( .D(n1459), .CP(clk), .Q(\memory[12][61] ) );
  CFD1QXL \memory_reg[12][60]  ( .D(n1460), .CP(clk), .Q(\memory[12][60] ) );
  CFD1QXL \memory_reg[12][59]  ( .D(n1461), .CP(clk), .Q(\memory[12][59] ) );
  CFD1QXL \memory_reg[12][58]  ( .D(n1462), .CP(clk), .Q(\memory[12][58] ) );
  CFD1QXL \memory_reg[12][57]  ( .D(n1463), .CP(clk), .Q(\memory[12][57] ) );
  CFD1QXL \memory_reg[12][56]  ( .D(n1464), .CP(clk), .Q(\memory[12][56] ) );
  CFD1QXL \memory_reg[12][55]  ( .D(n1465), .CP(clk), .Q(\memory[12][55] ) );
  CFD1QXL \memory_reg[12][54]  ( .D(n1466), .CP(clk), .Q(\memory[12][54] ) );
  CFD1QXL \memory_reg[12][53]  ( .D(n1467), .CP(clk), .Q(\memory[12][53] ) );
  CFD1QXL \memory_reg[12][52]  ( .D(n1468), .CP(clk), .Q(\memory[12][52] ) );
  CFD1QXL \memory_reg[12][51]  ( .D(n1469), .CP(clk), .Q(\memory[12][51] ) );
  CFD1QXL \memory_reg[12][50]  ( .D(n1470), .CP(clk), .Q(\memory[12][50] ) );
  CFD1QXL \memory_reg[12][49]  ( .D(n1471), .CP(clk), .Q(\memory[12][49] ) );
  CFD1QXL \memory_reg[12][48]  ( .D(n1472), .CP(clk), .Q(\memory[12][48] ) );
  CFD1QXL \memory_reg[12][47]  ( .D(n1473), .CP(clk), .Q(\memory[12][47] ) );
  CFD1QXL \memory_reg[12][46]  ( .D(n1474), .CP(clk), .Q(\memory[12][46] ) );
  CFD1QXL \memory_reg[12][45]  ( .D(n1475), .CP(clk), .Q(\memory[12][45] ) );
  CFD1QXL \memory_reg[12][44]  ( .D(n1476), .CP(clk), .Q(\memory[12][44] ) );
  CFD1QXL \memory_reg[12][43]  ( .D(n1477), .CP(clk), .Q(\memory[12][43] ) );
  CFD1QXL \memory_reg[12][42]  ( .D(n1478), .CP(clk), .Q(\memory[12][42] ) );
  CFD1QXL \memory_reg[12][41]  ( .D(n1479), .CP(clk), .Q(\memory[12][41] ) );
  CFD1QXL \memory_reg[12][40]  ( .D(n1480), .CP(clk), .Q(\memory[12][40] ) );
  CFD1QXL \memory_reg[12][39]  ( .D(n1481), .CP(clk), .Q(\memory[12][39] ) );
  CFD1QXL \memory_reg[12][38]  ( .D(n1482), .CP(clk), .Q(\memory[12][38] ) );
  CFD1QXL \memory_reg[12][37]  ( .D(n1483), .CP(clk), .Q(\memory[12][37] ) );
  CFD1QXL \memory_reg[12][36]  ( .D(n1484), .CP(clk), .Q(\memory[12][36] ) );
  CFD1QXL \memory_reg[12][35]  ( .D(n1485), .CP(clk), .Q(\memory[12][35] ) );
  CFD1QXL \memory_reg[12][34]  ( .D(n1486), .CP(clk), .Q(\memory[12][34] ) );
  CFD1QXL \memory_reg[12][33]  ( .D(n1487), .CP(clk), .Q(\memory[12][33] ) );
  CFD1QXL \memory_reg[12][32]  ( .D(n1488), .CP(clk), .Q(\memory[12][32] ) );
  CFD1QXL \memory_reg[12][31]  ( .D(n1489), .CP(clk), .Q(\memory[12][31] ) );
  CFD1QXL \memory_reg[12][30]  ( .D(n1490), .CP(clk), .Q(\memory[12][30] ) );
  CFD1QXL \memory_reg[12][29]  ( .D(n1491), .CP(clk), .Q(\memory[12][29] ) );
  CFD1QXL \memory_reg[12][28]  ( .D(n1492), .CP(clk), .Q(\memory[12][28] ) );
  CFD1QXL \memory_reg[12][27]  ( .D(n1493), .CP(clk), .Q(\memory[12][27] ) );
  CFD1QXL \memory_reg[12][26]  ( .D(n1494), .CP(clk), .Q(\memory[12][26] ) );
  CFD1QXL \memory_reg[12][25]  ( .D(n1495), .CP(clk), .Q(\memory[12][25] ) );
  CFD1QXL \memory_reg[12][24]  ( .D(n1496), .CP(clk), .Q(\memory[12][24] ) );
  CFD1QXL \memory_reg[12][23]  ( .D(n1497), .CP(clk), .Q(\memory[12][23] ) );
  CFD1QXL \memory_reg[12][22]  ( .D(n1498), .CP(clk), .Q(\memory[12][22] ) );
  CFD1QXL \memory_reg[12][21]  ( .D(n1499), .CP(clk), .Q(\memory[12][21] ) );
  CFD1QXL \memory_reg[12][20]  ( .D(n1500), .CP(clk), .Q(\memory[12][20] ) );
  CFD1QXL \memory_reg[12][19]  ( .D(n1501), .CP(clk), .Q(\memory[12][19] ) );
  CFD1QXL \memory_reg[12][18]  ( .D(n1502), .CP(clk), .Q(\memory[12][18] ) );
  CFD1QXL \memory_reg[12][17]  ( .D(n1503), .CP(clk), .Q(\memory[12][17] ) );
  CFD1QXL \memory_reg[12][16]  ( .D(n1504), .CP(clk), .Q(\memory[12][16] ) );
  CFD1QXL \memory_reg[12][15]  ( .D(n1505), .CP(clk), .Q(\memory[12][15] ) );
  CFD1QXL \memory_reg[12][14]  ( .D(n1506), .CP(clk), .Q(\memory[12][14] ) );
  CFD1QXL \memory_reg[12][13]  ( .D(n1507), .CP(clk), .Q(\memory[12][13] ) );
  CFD1QXL \memory_reg[12][12]  ( .D(n1508), .CP(clk), .Q(\memory[12][12] ) );
  CFD1QXL \memory_reg[12][11]  ( .D(n1509), .CP(clk), .Q(\memory[12][11] ) );
  CFD1QXL \memory_reg[12][10]  ( .D(n1510), .CP(clk), .Q(\memory[12][10] ) );
  CFD1QXL \memory_reg[12][9]  ( .D(n1511), .CP(clk), .Q(\memory[12][9] ) );
  CFD1QXL \memory_reg[12][8]  ( .D(n1512), .CP(clk), .Q(\memory[12][8] ) );
  CFD1QXL \memory_reg[12][7]  ( .D(n1513), .CP(clk), .Q(\memory[12][7] ) );
  CFD1QXL \memory_reg[12][6]  ( .D(n1514), .CP(clk), .Q(\memory[12][6] ) );
  CFD1QXL \memory_reg[12][5]  ( .D(n1515), .CP(clk), .Q(\memory[12][5] ) );
  CFD1QXL \memory_reg[12][4]  ( .D(n1516), .CP(clk), .Q(\memory[12][4] ) );
  CFD1QXL \memory_reg[12][3]  ( .D(n1517), .CP(clk), .Q(\memory[12][3] ) );
  CFD1QXL \memory_reg[12][2]  ( .D(n1518), .CP(clk), .Q(\memory[12][2] ) );
  CFD1QXL \memory_reg[12][1]  ( .D(n1519), .CP(clk), .Q(\memory[12][1] ) );
  CFD1QXL \memory_reg[12][0]  ( .D(n1520), .CP(clk), .Q(\memory[12][0] ) );
  CFD1QXL \memory_reg[11][63]  ( .D(n1528), .CP(clk), .Q(\memory[11][63] ) );
  CFD1QXL \memory_reg[11][62]  ( .D(n1529), .CP(clk), .Q(\memory[11][62] ) );
  CFD1QXL \memory_reg[11][61]  ( .D(n1530), .CP(clk), .Q(\memory[11][61] ) );
  CFD1QXL \memory_reg[11][60]  ( .D(n1531), .CP(clk), .Q(\memory[11][60] ) );
  CFD1QXL \memory_reg[11][59]  ( .D(n1532), .CP(clk), .Q(\memory[11][59] ) );
  CFD1QXL \memory_reg[11][58]  ( .D(n1533), .CP(clk), .Q(\memory[11][58] ) );
  CFD1QXL \memory_reg[11][57]  ( .D(n1534), .CP(clk), .Q(\memory[11][57] ) );
  CFD1QXL \memory_reg[11][56]  ( .D(n1535), .CP(clk), .Q(\memory[11][56] ) );
  CFD1QXL \memory_reg[11][55]  ( .D(n1536), .CP(clk), .Q(\memory[11][55] ) );
  CFD1QXL \memory_reg[11][54]  ( .D(n1537), .CP(clk), .Q(\memory[11][54] ) );
  CFD1QXL \memory_reg[11][53]  ( .D(n1538), .CP(clk), .Q(\memory[11][53] ) );
  CFD1QXL \memory_reg[11][52]  ( .D(n1539), .CP(clk), .Q(\memory[11][52] ) );
  CFD1QXL \memory_reg[11][51]  ( .D(n1540), .CP(clk), .Q(\memory[11][51] ) );
  CFD1QXL \memory_reg[11][50]  ( .D(n1541), .CP(clk), .Q(\memory[11][50] ) );
  CFD1QXL \memory_reg[11][49]  ( .D(n1542), .CP(clk), .Q(\memory[11][49] ) );
  CFD1QXL \memory_reg[11][48]  ( .D(n1543), .CP(clk), .Q(\memory[11][48] ) );
  CFD1QXL \memory_reg[11][47]  ( .D(n1544), .CP(clk), .Q(\memory[11][47] ) );
  CFD1QXL \memory_reg[11][46]  ( .D(n1545), .CP(clk), .Q(\memory[11][46] ) );
  CFD1QXL \memory_reg[11][45]  ( .D(n1546), .CP(clk), .Q(\memory[11][45] ) );
  CFD1QXL \memory_reg[11][44]  ( .D(n1547), .CP(clk), .Q(\memory[11][44] ) );
  CFD1QXL \memory_reg[11][43]  ( .D(n1548), .CP(clk), .Q(\memory[11][43] ) );
  CFD1QXL \memory_reg[11][42]  ( .D(n1549), .CP(clk), .Q(\memory[11][42] ) );
  CFD1QXL \memory_reg[11][41]  ( .D(n1550), .CP(clk), .Q(\memory[11][41] ) );
  CFD1QXL \memory_reg[11][40]  ( .D(n1551), .CP(clk), .Q(\memory[11][40] ) );
  CFD1QXL \memory_reg[11][39]  ( .D(n1552), .CP(clk), .Q(\memory[11][39] ) );
  CFD1QXL \memory_reg[11][38]  ( .D(n1553), .CP(clk), .Q(\memory[11][38] ) );
  CFD1QXL \memory_reg[11][37]  ( .D(n1554), .CP(clk), .Q(\memory[11][37] ) );
  CFD1QXL \memory_reg[11][36]  ( .D(n1555), .CP(clk), .Q(\memory[11][36] ) );
  CFD1QXL \memory_reg[11][35]  ( .D(n1556), .CP(clk), .Q(\memory[11][35] ) );
  CFD1QXL \memory_reg[11][34]  ( .D(n1557), .CP(clk), .Q(\memory[11][34] ) );
  CFD1QXL \memory_reg[11][33]  ( .D(n1558), .CP(clk), .Q(\memory[11][33] ) );
  CFD1QXL \memory_reg[11][32]  ( .D(n1559), .CP(clk), .Q(\memory[11][32] ) );
  CFD1QXL \memory_reg[11][31]  ( .D(n1560), .CP(clk), .Q(\memory[11][31] ) );
  CFD1QXL \memory_reg[11][30]  ( .D(n1561), .CP(clk), .Q(\memory[11][30] ) );
  CFD1QXL \memory_reg[11][29]  ( .D(n1562), .CP(clk), .Q(\memory[11][29] ) );
  CFD1QXL \memory_reg[11][28]  ( .D(n1563), .CP(clk), .Q(\memory[11][28] ) );
  CFD1QXL \memory_reg[11][27]  ( .D(n1564), .CP(clk), .Q(\memory[11][27] ) );
  CFD1QXL \memory_reg[11][26]  ( .D(n1565), .CP(clk), .Q(\memory[11][26] ) );
  CFD1QXL \memory_reg[11][25]  ( .D(n1566), .CP(clk), .Q(\memory[11][25] ) );
  CFD1QXL \memory_reg[11][24]  ( .D(n1567), .CP(clk), .Q(\memory[11][24] ) );
  CFD1QXL \memory_reg[11][23]  ( .D(n1568), .CP(clk), .Q(\memory[11][23] ) );
  CFD1QXL \memory_reg[11][22]  ( .D(n1569), .CP(clk), .Q(\memory[11][22] ) );
  CFD1QXL \memory_reg[11][21]  ( .D(n1570), .CP(clk), .Q(\memory[11][21] ) );
  CFD1QXL \memory_reg[11][20]  ( .D(n1571), .CP(clk), .Q(\memory[11][20] ) );
  CFD1QXL \memory_reg[11][19]  ( .D(n1572), .CP(clk), .Q(\memory[11][19] ) );
  CFD1QXL \memory_reg[11][18]  ( .D(n1573), .CP(clk), .Q(\memory[11][18] ) );
  CFD1QXL \memory_reg[11][17]  ( .D(n1574), .CP(clk), .Q(\memory[11][17] ) );
  CFD1QXL \memory_reg[11][16]  ( .D(n1575), .CP(clk), .Q(\memory[11][16] ) );
  CFD1QXL \memory_reg[11][15]  ( .D(n1576), .CP(clk), .Q(\memory[11][15] ) );
  CFD1QXL \memory_reg[11][14]  ( .D(n1577), .CP(clk), .Q(\memory[11][14] ) );
  CFD1QXL \memory_reg[11][13]  ( .D(n1578), .CP(clk), .Q(\memory[11][13] ) );
  CFD1QXL \memory_reg[11][12]  ( .D(n1579), .CP(clk), .Q(\memory[11][12] ) );
  CFD1QXL \memory_reg[11][11]  ( .D(n1580), .CP(clk), .Q(\memory[11][11] ) );
  CFD1QXL \memory_reg[11][10]  ( .D(n1581), .CP(clk), .Q(\memory[11][10] ) );
  CFD1QXL \memory_reg[11][9]  ( .D(n1582), .CP(clk), .Q(\memory[11][9] ) );
  CFD1QXL \memory_reg[11][8]  ( .D(n1583), .CP(clk), .Q(\memory[11][8] ) );
  CFD1QXL \memory_reg[11][7]  ( .D(n1584), .CP(clk), .Q(\memory[11][7] ) );
  CFD1QXL \memory_reg[11][6]  ( .D(n1585), .CP(clk), .Q(\memory[11][6] ) );
  CFD1QXL \memory_reg[11][5]  ( .D(n1586), .CP(clk), .Q(\memory[11][5] ) );
  CFD1QXL \memory_reg[11][4]  ( .D(n1587), .CP(clk), .Q(\memory[11][4] ) );
  CFD1QXL \memory_reg[11][3]  ( .D(n1588), .CP(clk), .Q(\memory[11][3] ) );
  CFD1QXL \memory_reg[11][2]  ( .D(n1589), .CP(clk), .Q(\memory[11][2] ) );
  CFD1QXL \memory_reg[11][1]  ( .D(n1590), .CP(clk), .Q(\memory[11][1] ) );
  CFD1QXL \memory_reg[11][0]  ( .D(n1591), .CP(clk), .Q(\memory[11][0] ) );
  CFD1QXL \memory_reg[10][63]  ( .D(n1599), .CP(clk), .Q(\memory[10][63] ) );
  CFD1QXL \memory_reg[10][62]  ( .D(n1600), .CP(clk), .Q(\memory[10][62] ) );
  CFD1QXL \memory_reg[10][61]  ( .D(n1601), .CP(clk), .Q(\memory[10][61] ) );
  CFD1QXL \memory_reg[10][60]  ( .D(n1602), .CP(clk), .Q(\memory[10][60] ) );
  CFD1QXL \memory_reg[10][59]  ( .D(n1603), .CP(clk), .Q(\memory[10][59] ) );
  CFD1QXL \memory_reg[10][58]  ( .D(n1604), .CP(clk), .Q(\memory[10][58] ) );
  CFD1QXL \memory_reg[10][57]  ( .D(n1605), .CP(clk), .Q(\memory[10][57] ) );
  CFD1QXL \memory_reg[10][56]  ( .D(n1606), .CP(clk), .Q(\memory[10][56] ) );
  CFD1QXL \memory_reg[10][55]  ( .D(n1607), .CP(clk), .Q(\memory[10][55] ) );
  CFD1QXL \memory_reg[10][54]  ( .D(n1608), .CP(clk), .Q(\memory[10][54] ) );
  CFD1QXL \memory_reg[10][53]  ( .D(n1609), .CP(clk), .Q(\memory[10][53] ) );
  CFD1QXL \memory_reg[10][52]  ( .D(n1610), .CP(clk), .Q(\memory[10][52] ) );
  CFD1QXL \memory_reg[10][51]  ( .D(n1611), .CP(clk), .Q(\memory[10][51] ) );
  CFD1QXL \memory_reg[10][50]  ( .D(n1612), .CP(clk), .Q(\memory[10][50] ) );
  CFD1QXL \memory_reg[10][49]  ( .D(n1613), .CP(clk), .Q(\memory[10][49] ) );
  CFD1QXL \memory_reg[10][48]  ( .D(n1614), .CP(clk), .Q(\memory[10][48] ) );
  CFD1QXL \memory_reg[10][47]  ( .D(n1615), .CP(clk), .Q(\memory[10][47] ) );
  CFD1QXL \memory_reg[10][46]  ( .D(n1616), .CP(clk), .Q(\memory[10][46] ) );
  CFD1QXL \memory_reg[10][45]  ( .D(n1617), .CP(clk), .Q(\memory[10][45] ) );
  CFD1QXL \memory_reg[10][44]  ( .D(n1618), .CP(clk), .Q(\memory[10][44] ) );
  CFD1QXL \memory_reg[10][43]  ( .D(n1619), .CP(clk), .Q(\memory[10][43] ) );
  CFD1QXL \memory_reg[10][42]  ( .D(n1620), .CP(clk), .Q(\memory[10][42] ) );
  CFD1QXL \memory_reg[10][41]  ( .D(n1621), .CP(clk), .Q(\memory[10][41] ) );
  CFD1QXL \memory_reg[10][40]  ( .D(n1622), .CP(clk), .Q(\memory[10][40] ) );
  CFD1QXL \memory_reg[10][39]  ( .D(n1623), .CP(clk), .Q(\memory[10][39] ) );
  CFD1QXL \memory_reg[10][38]  ( .D(n1624), .CP(clk), .Q(\memory[10][38] ) );
  CFD1QXL \memory_reg[10][37]  ( .D(n1625), .CP(clk), .Q(\memory[10][37] ) );
  CFD1QXL \memory_reg[10][36]  ( .D(n1626), .CP(clk), .Q(\memory[10][36] ) );
  CFD1QXL \memory_reg[10][35]  ( .D(n1627), .CP(clk), .Q(\memory[10][35] ) );
  CFD1QXL \memory_reg[10][34]  ( .D(n1628), .CP(clk), .Q(\memory[10][34] ) );
  CFD1QXL \memory_reg[10][33]  ( .D(n1629), .CP(clk), .Q(\memory[10][33] ) );
  CFD1QXL \memory_reg[10][32]  ( .D(n1630), .CP(clk), .Q(\memory[10][32] ) );
  CFD1QXL \memory_reg[10][31]  ( .D(n1631), .CP(clk), .Q(\memory[10][31] ) );
  CFD1QXL \memory_reg[10][30]  ( .D(n1632), .CP(clk), .Q(\memory[10][30] ) );
  CFD1QXL \memory_reg[10][29]  ( .D(n1633), .CP(clk), .Q(\memory[10][29] ) );
  CFD1QXL \memory_reg[10][28]  ( .D(n1634), .CP(clk), .Q(\memory[10][28] ) );
  CFD1QXL \memory_reg[10][27]  ( .D(n1635), .CP(clk), .Q(\memory[10][27] ) );
  CFD1QXL \memory_reg[10][26]  ( .D(n1636), .CP(clk), .Q(\memory[10][26] ) );
  CFD1QXL \memory_reg[10][25]  ( .D(n1637), .CP(clk), .Q(\memory[10][25] ) );
  CFD1QXL \memory_reg[10][24]  ( .D(n1638), .CP(clk), .Q(\memory[10][24] ) );
  CFD1QXL \memory_reg[10][23]  ( .D(n1639), .CP(clk), .Q(\memory[10][23] ) );
  CFD1QXL \memory_reg[10][22]  ( .D(n1640), .CP(clk), .Q(\memory[10][22] ) );
  CFD1QXL \memory_reg[10][21]  ( .D(n1641), .CP(clk), .Q(\memory[10][21] ) );
  CFD1QXL \memory_reg[10][20]  ( .D(n1642), .CP(clk), .Q(\memory[10][20] ) );
  CFD1QXL \memory_reg[10][19]  ( .D(n1643), .CP(clk), .Q(\memory[10][19] ) );
  CFD1QXL \memory_reg[10][18]  ( .D(n1644), .CP(clk), .Q(\memory[10][18] ) );
  CFD1QXL \memory_reg[10][17]  ( .D(n1645), .CP(clk), .Q(\memory[10][17] ) );
  CFD1QXL \memory_reg[10][16]  ( .D(n1646), .CP(clk), .Q(\memory[10][16] ) );
  CFD1QXL \memory_reg[10][15]  ( .D(n1647), .CP(clk), .Q(\memory[10][15] ) );
  CFD1QXL \memory_reg[10][14]  ( .D(n1648), .CP(clk), .Q(\memory[10][14] ) );
  CFD1QXL \memory_reg[10][13]  ( .D(n1649), .CP(clk), .Q(\memory[10][13] ) );
  CFD1QXL \memory_reg[10][12]  ( .D(n1650), .CP(clk), .Q(\memory[10][12] ) );
  CFD1QXL \memory_reg[10][11]  ( .D(n1651), .CP(clk), .Q(\memory[10][11] ) );
  CFD1QXL \memory_reg[10][10]  ( .D(n1652), .CP(clk), .Q(\memory[10][10] ) );
  CFD1QXL \memory_reg[10][9]  ( .D(n1653), .CP(clk), .Q(\memory[10][9] ) );
  CFD1QXL \memory_reg[10][8]  ( .D(n1654), .CP(clk), .Q(\memory[10][8] ) );
  CFD1QXL \memory_reg[10][7]  ( .D(n1655), .CP(clk), .Q(\memory[10][7] ) );
  CFD1QXL \memory_reg[10][6]  ( .D(n1656), .CP(clk), .Q(\memory[10][6] ) );
  CFD1QXL \memory_reg[10][5]  ( .D(n1657), .CP(clk), .Q(\memory[10][5] ) );
  CFD1QXL \memory_reg[10][4]  ( .D(n1658), .CP(clk), .Q(\memory[10][4] ) );
  CFD1QXL \memory_reg[10][3]  ( .D(n1659), .CP(clk), .Q(\memory[10][3] ) );
  CFD1QXL \memory_reg[10][2]  ( .D(n1660), .CP(clk), .Q(\memory[10][2] ) );
  CFD1QXL \memory_reg[10][1]  ( .D(n1661), .CP(clk), .Q(\memory[10][1] ) );
  CFD1QXL \memory_reg[10][0]  ( .D(n1662), .CP(clk), .Q(\memory[10][0] ) );
  CFD1QXL \memory_reg[9][63]  ( .D(n1670), .CP(clk), .Q(\memory[9][63] ) );
  CFD1QXL \memory_reg[9][62]  ( .D(n1671), .CP(clk), .Q(\memory[9][62] ) );
  CFD1QXL \memory_reg[9][61]  ( .D(n1672), .CP(clk), .Q(\memory[9][61] ) );
  CFD1QXL \memory_reg[9][60]  ( .D(n1673), .CP(clk), .Q(\memory[9][60] ) );
  CFD1QXL \memory_reg[9][59]  ( .D(n1674), .CP(clk), .Q(\memory[9][59] ) );
  CFD1QXL \memory_reg[9][58]  ( .D(n1675), .CP(clk), .Q(\memory[9][58] ) );
  CFD1QXL \memory_reg[9][57]  ( .D(n1676), .CP(clk), .Q(\memory[9][57] ) );
  CFD1QXL \memory_reg[9][56]  ( .D(n1677), .CP(clk), .Q(\memory[9][56] ) );
  CFD1QXL \memory_reg[9][55]  ( .D(n1678), .CP(clk), .Q(\memory[9][55] ) );
  CFD1QXL \memory_reg[9][54]  ( .D(n1679), .CP(clk), .Q(\memory[9][54] ) );
  CFD1QXL \memory_reg[9][53]  ( .D(n1680), .CP(clk), .Q(\memory[9][53] ) );
  CFD1QXL \memory_reg[9][52]  ( .D(n1681), .CP(clk), .Q(\memory[9][52] ) );
  CFD1QXL \memory_reg[9][51]  ( .D(n1682), .CP(clk), .Q(\memory[9][51] ) );
  CFD1QXL \memory_reg[9][50]  ( .D(n1683), .CP(clk), .Q(\memory[9][50] ) );
  CFD1QXL \memory_reg[9][49]  ( .D(n1684), .CP(clk), .Q(\memory[9][49] ) );
  CFD1QXL \memory_reg[9][48]  ( .D(n1685), .CP(clk), .Q(\memory[9][48] ) );
  CFD1QXL \memory_reg[9][47]  ( .D(n1686), .CP(clk), .Q(\memory[9][47] ) );
  CFD1QXL \memory_reg[9][46]  ( .D(n1687), .CP(clk), .Q(\memory[9][46] ) );
  CFD1QXL \memory_reg[9][45]  ( .D(n1688), .CP(clk), .Q(\memory[9][45] ) );
  CFD1QXL \memory_reg[9][44]  ( .D(n1689), .CP(clk), .Q(\memory[9][44] ) );
  CFD1QXL \memory_reg[9][43]  ( .D(n1690), .CP(clk), .Q(\memory[9][43] ) );
  CFD1QXL \memory_reg[9][42]  ( .D(n1691), .CP(clk), .Q(\memory[9][42] ) );
  CFD1QXL \memory_reg[9][41]  ( .D(n1692), .CP(clk), .Q(\memory[9][41] ) );
  CFD1QXL \memory_reg[9][40]  ( .D(n1693), .CP(clk), .Q(\memory[9][40] ) );
  CFD1QXL \memory_reg[9][39]  ( .D(n1694), .CP(clk), .Q(\memory[9][39] ) );
  CFD1QXL \memory_reg[9][38]  ( .D(n1695), .CP(clk), .Q(\memory[9][38] ) );
  CFD1QXL \memory_reg[9][37]  ( .D(n1696), .CP(clk), .Q(\memory[9][37] ) );
  CFD1QXL \memory_reg[9][36]  ( .D(n1697), .CP(clk), .Q(\memory[9][36] ) );
  CFD1QXL \memory_reg[9][35]  ( .D(n1698), .CP(clk), .Q(\memory[9][35] ) );
  CFD1QXL \memory_reg[9][34]  ( .D(n1699), .CP(clk), .Q(\memory[9][34] ) );
  CFD1QXL \memory_reg[9][33]  ( .D(n1700), .CP(clk), .Q(\memory[9][33] ) );
  CFD1QXL \memory_reg[9][32]  ( .D(n1701), .CP(clk), .Q(\memory[9][32] ) );
  CFD1QXL \memory_reg[9][31]  ( .D(n1702), .CP(clk), .Q(\memory[9][31] ) );
  CFD1QXL \memory_reg[9][30]  ( .D(n1703), .CP(clk), .Q(\memory[9][30] ) );
  CFD1QXL \memory_reg[9][29]  ( .D(n1704), .CP(clk), .Q(\memory[9][29] ) );
  CFD1QXL \memory_reg[9][28]  ( .D(n1705), .CP(clk), .Q(\memory[9][28] ) );
  CFD1QXL \memory_reg[9][27]  ( .D(n1706), .CP(clk), .Q(\memory[9][27] ) );
  CFD1QXL \memory_reg[9][26]  ( .D(n1707), .CP(clk), .Q(\memory[9][26] ) );
  CFD1QXL \memory_reg[9][25]  ( .D(n1708), .CP(clk), .Q(\memory[9][25] ) );
  CFD1QXL \memory_reg[9][24]  ( .D(n1709), .CP(clk), .Q(\memory[9][24] ) );
  CFD1QXL \memory_reg[9][23]  ( .D(n1710), .CP(clk), .Q(\memory[9][23] ) );
  CFD1QXL \memory_reg[9][22]  ( .D(n1711), .CP(clk), .Q(\memory[9][22] ) );
  CFD1QXL \memory_reg[9][21]  ( .D(n1712), .CP(clk), .Q(\memory[9][21] ) );
  CFD1QXL \memory_reg[9][20]  ( .D(n1713), .CP(clk), .Q(\memory[9][20] ) );
  CFD1QXL \memory_reg[9][19]  ( .D(n1714), .CP(clk), .Q(\memory[9][19] ) );
  CFD1QXL \memory_reg[9][18]  ( .D(n1715), .CP(clk), .Q(\memory[9][18] ) );
  CFD1QXL \memory_reg[9][17]  ( .D(n1716), .CP(clk), .Q(\memory[9][17] ) );
  CFD1QXL \memory_reg[9][16]  ( .D(n1717), .CP(clk), .Q(\memory[9][16] ) );
  CFD1QXL \memory_reg[9][15]  ( .D(n1718), .CP(clk), .Q(\memory[9][15] ) );
  CFD1QXL \memory_reg[9][14]  ( .D(n1719), .CP(clk), .Q(\memory[9][14] ) );
  CFD1QXL \memory_reg[9][13]  ( .D(n1720), .CP(clk), .Q(\memory[9][13] ) );
  CFD1QXL \memory_reg[9][12]  ( .D(n1721), .CP(clk), .Q(\memory[9][12] ) );
  CFD1QXL \memory_reg[9][11]  ( .D(n1722), .CP(clk), .Q(\memory[9][11] ) );
  CFD1QXL \memory_reg[9][10]  ( .D(n1723), .CP(clk), .Q(\memory[9][10] ) );
  CFD1QXL \memory_reg[9][9]  ( .D(n1724), .CP(clk), .Q(\memory[9][9] ) );
  CFD1QXL \memory_reg[9][8]  ( .D(n1725), .CP(clk), .Q(\memory[9][8] ) );
  CFD1QXL \memory_reg[9][7]  ( .D(n1726), .CP(clk), .Q(\memory[9][7] ) );
  CFD1QXL \memory_reg[9][6]  ( .D(n1727), .CP(clk), .Q(\memory[9][6] ) );
  CFD1QXL \memory_reg[9][5]  ( .D(n1728), .CP(clk), .Q(\memory[9][5] ) );
  CFD1QXL \memory_reg[9][4]  ( .D(n1729), .CP(clk), .Q(\memory[9][4] ) );
  CFD1QXL \memory_reg[9][3]  ( .D(n1730), .CP(clk), .Q(\memory[9][3] ) );
  CFD1QXL \memory_reg[9][2]  ( .D(n1731), .CP(clk), .Q(\memory[9][2] ) );
  CFD1QXL \memory_reg[9][1]  ( .D(n1732), .CP(clk), .Q(\memory[9][1] ) );
  CFD1QXL \memory_reg[9][0]  ( .D(n1733), .CP(clk), .Q(\memory[9][0] ) );
  CFD1QXL \memory_reg[8][63]  ( .D(n1741), .CP(clk), .Q(\memory[8][63] ) );
  CFD1QXL \memory_reg[8][62]  ( .D(n1742), .CP(clk), .Q(\memory[8][62] ) );
  CFD1QXL \memory_reg[8][61]  ( .D(n1743), .CP(clk), .Q(\memory[8][61] ) );
  CFD1QXL \memory_reg[8][60]  ( .D(n1744), .CP(clk), .Q(\memory[8][60] ) );
  CFD1QXL \memory_reg[8][59]  ( .D(n1745), .CP(clk), .Q(\memory[8][59] ) );
  CFD1QXL \memory_reg[8][58]  ( .D(n1746), .CP(clk), .Q(\memory[8][58] ) );
  CFD1QXL \memory_reg[8][57]  ( .D(n1747), .CP(clk), .Q(\memory[8][57] ) );
  CFD1QXL \memory_reg[8][56]  ( .D(n1748), .CP(clk), .Q(\memory[8][56] ) );
  CFD1QXL \memory_reg[8][55]  ( .D(n1749), .CP(clk), .Q(\memory[8][55] ) );
  CFD1QXL \memory_reg[8][54]  ( .D(n1750), .CP(clk), .Q(\memory[8][54] ) );
  CFD1QXL \memory_reg[8][53]  ( .D(n1751), .CP(clk), .Q(\memory[8][53] ) );
  CFD1QXL \memory_reg[8][52]  ( .D(n1752), .CP(clk), .Q(\memory[8][52] ) );
  CFD1QXL \memory_reg[8][51]  ( .D(n1753), .CP(clk), .Q(\memory[8][51] ) );
  CFD1QXL \memory_reg[8][50]  ( .D(n1754), .CP(clk), .Q(\memory[8][50] ) );
  CFD1QXL \memory_reg[8][49]  ( .D(n1755), .CP(clk), .Q(\memory[8][49] ) );
  CFD1QXL \memory_reg[8][48]  ( .D(n1756), .CP(clk), .Q(\memory[8][48] ) );
  CFD1QXL \memory_reg[8][47]  ( .D(n1757), .CP(clk), .Q(\memory[8][47] ) );
  CFD1QXL \memory_reg[8][46]  ( .D(n1758), .CP(clk), .Q(\memory[8][46] ) );
  CFD1QXL \memory_reg[8][45]  ( .D(n1759), .CP(clk), .Q(\memory[8][45] ) );
  CFD1QXL \memory_reg[8][44]  ( .D(n1760), .CP(clk), .Q(\memory[8][44] ) );
  CFD1QXL \memory_reg[8][43]  ( .D(n1761), .CP(clk), .Q(\memory[8][43] ) );
  CFD1QXL \memory_reg[8][42]  ( .D(n1762), .CP(clk), .Q(\memory[8][42] ) );
  CFD1QXL \memory_reg[8][41]  ( .D(n1763), .CP(clk), .Q(\memory[8][41] ) );
  CFD1QXL \memory_reg[8][40]  ( .D(n1764), .CP(clk), .Q(\memory[8][40] ) );
  CFD1QXL \memory_reg[8][39]  ( .D(n1765), .CP(clk), .Q(\memory[8][39] ) );
  CFD1QXL \memory_reg[8][38]  ( .D(n1766), .CP(clk), .Q(\memory[8][38] ) );
  CFD1QXL \memory_reg[8][37]  ( .D(n1767), .CP(clk), .Q(\memory[8][37] ) );
  CFD1QXL \memory_reg[8][36]  ( .D(n1768), .CP(clk), .Q(\memory[8][36] ) );
  CFD1QXL \memory_reg[8][35]  ( .D(n1769), .CP(clk), .Q(\memory[8][35] ) );
  CFD1QXL \memory_reg[8][34]  ( .D(n1770), .CP(clk), .Q(\memory[8][34] ) );
  CFD1QXL \memory_reg[8][33]  ( .D(n1771), .CP(clk), .Q(\memory[8][33] ) );
  CFD1QXL \memory_reg[8][32]  ( .D(n1772), .CP(clk), .Q(\memory[8][32] ) );
  CFD1QXL \memory_reg[8][31]  ( .D(n1773), .CP(clk), .Q(\memory[8][31] ) );
  CFD1QXL \memory_reg[8][30]  ( .D(n1774), .CP(clk), .Q(\memory[8][30] ) );
  CFD1QXL \memory_reg[8][29]  ( .D(n1775), .CP(clk), .Q(\memory[8][29] ) );
  CFD1QXL \memory_reg[8][28]  ( .D(n1776), .CP(clk), .Q(\memory[8][28] ) );
  CFD1QXL \memory_reg[8][27]  ( .D(n1777), .CP(clk), .Q(\memory[8][27] ) );
  CFD1QXL \memory_reg[8][26]  ( .D(n1778), .CP(clk), .Q(\memory[8][26] ) );
  CFD1QXL \memory_reg[8][25]  ( .D(n1779), .CP(clk), .Q(\memory[8][25] ) );
  CFD1QXL \memory_reg[8][24]  ( .D(n1780), .CP(clk), .Q(\memory[8][24] ) );
  CFD1QXL \memory_reg[8][23]  ( .D(n1781), .CP(clk), .Q(\memory[8][23] ) );
  CFD1QXL \memory_reg[8][22]  ( .D(n1782), .CP(clk), .Q(\memory[8][22] ) );
  CFD1QXL \memory_reg[8][21]  ( .D(n1783), .CP(clk), .Q(\memory[8][21] ) );
  CFD1QXL \memory_reg[8][20]  ( .D(n1784), .CP(clk), .Q(\memory[8][20] ) );
  CFD1QXL \memory_reg[8][19]  ( .D(n1785), .CP(clk), .Q(\memory[8][19] ) );
  CFD1QXL \memory_reg[8][18]  ( .D(n1786), .CP(clk), .Q(\memory[8][18] ) );
  CFD1QXL \memory_reg[8][17]  ( .D(n1787), .CP(clk), .Q(\memory[8][17] ) );
  CFD1QXL \memory_reg[8][16]  ( .D(n1788), .CP(clk), .Q(\memory[8][16] ) );
  CFD1QXL \memory_reg[8][15]  ( .D(n1789), .CP(clk), .Q(\memory[8][15] ) );
  CFD1QXL \memory_reg[8][14]  ( .D(n1790), .CP(clk), .Q(\memory[8][14] ) );
  CFD1QXL \memory_reg[8][13]  ( .D(n1791), .CP(clk), .Q(\memory[8][13] ) );
  CFD1QXL \memory_reg[8][12]  ( .D(n1792), .CP(clk), .Q(\memory[8][12] ) );
  CFD1QXL \memory_reg[8][11]  ( .D(n1793), .CP(clk), .Q(\memory[8][11] ) );
  CFD1QXL \memory_reg[8][10]  ( .D(n1794), .CP(clk), .Q(\memory[8][10] ) );
  CFD1QXL \memory_reg[8][9]  ( .D(n1795), .CP(clk), .Q(\memory[8][9] ) );
  CFD1QXL \memory_reg[8][8]  ( .D(n1796), .CP(clk), .Q(\memory[8][8] ) );
  CFD1QXL \memory_reg[8][7]  ( .D(n1797), .CP(clk), .Q(\memory[8][7] ) );
  CFD1QXL \memory_reg[8][6]  ( .D(n1798), .CP(clk), .Q(\memory[8][6] ) );
  CFD1QXL \memory_reg[8][5]  ( .D(n1799), .CP(clk), .Q(\memory[8][5] ) );
  CFD1QXL \memory_reg[8][4]  ( .D(n1800), .CP(clk), .Q(\memory[8][4] ) );
  CFD1QXL \memory_reg[8][3]  ( .D(n1801), .CP(clk), .Q(\memory[8][3] ) );
  CFD1QXL \memory_reg[8][2]  ( .D(n1802), .CP(clk), .Q(\memory[8][2] ) );
  CFD1QXL \memory_reg[8][1]  ( .D(n1803), .CP(clk), .Q(\memory[8][1] ) );
  CFD1QXL \memory_reg[8][0]  ( .D(n1804), .CP(clk), .Q(\memory[8][0] ) );
  CFD1QXL \memory_reg[6][63]  ( .D(n1883), .CP(clk), .Q(\memory[6][63] ) );
  CFD1QXL \memory_reg[6][62]  ( .D(n1884), .CP(clk), .Q(\memory[6][62] ) );
  CFD1QXL \memory_reg[6][61]  ( .D(n1885), .CP(clk), .Q(\memory[6][61] ) );
  CFD1QXL \memory_reg[6][60]  ( .D(n1886), .CP(clk), .Q(\memory[6][60] ) );
  CFD1QXL \memory_reg[6][59]  ( .D(n1887), .CP(clk), .Q(\memory[6][59] ) );
  CFD1QXL \memory_reg[6][58]  ( .D(n1888), .CP(clk), .Q(\memory[6][58] ) );
  CFD1QXL \memory_reg[6][57]  ( .D(n1889), .CP(clk), .Q(\memory[6][57] ) );
  CFD1QXL \memory_reg[6][56]  ( .D(n1890), .CP(clk), .Q(\memory[6][56] ) );
  CFD1QXL \memory_reg[6][55]  ( .D(n1891), .CP(clk), .Q(\memory[6][55] ) );
  CFD1QXL \memory_reg[6][54]  ( .D(n1892), .CP(clk), .Q(\memory[6][54] ) );
  CFD1QXL \memory_reg[6][53]  ( .D(n1893), .CP(clk), .Q(\memory[6][53] ) );
  CFD1QXL \memory_reg[6][52]  ( .D(n1894), .CP(clk), .Q(\memory[6][52] ) );
  CFD1QXL \memory_reg[6][51]  ( .D(n1895), .CP(clk), .Q(\memory[6][51] ) );
  CFD1QXL \memory_reg[6][50]  ( .D(n1896), .CP(clk), .Q(\memory[6][50] ) );
  CFD1QXL \memory_reg[6][49]  ( .D(n1897), .CP(clk), .Q(\memory[6][49] ) );
  CFD1QXL \memory_reg[6][48]  ( .D(n1898), .CP(clk), .Q(\memory[6][48] ) );
  CFD1QXL \memory_reg[6][47]  ( .D(n1899), .CP(clk), .Q(\memory[6][47] ) );
  CFD1QXL \memory_reg[6][46]  ( .D(n1900), .CP(clk), .Q(\memory[6][46] ) );
  CFD1QXL \memory_reg[6][45]  ( .D(n1901), .CP(clk), .Q(\memory[6][45] ) );
  CFD1QXL \memory_reg[6][44]  ( .D(n1902), .CP(clk), .Q(\memory[6][44] ) );
  CFD1QXL \memory_reg[6][43]  ( .D(n1903), .CP(clk), .Q(\memory[6][43] ) );
  CFD1QXL \memory_reg[6][42]  ( .D(n1904), .CP(clk), .Q(\memory[6][42] ) );
  CFD1QXL \memory_reg[6][41]  ( .D(n1905), .CP(clk), .Q(\memory[6][41] ) );
  CFD1QXL \memory_reg[6][40]  ( .D(n1906), .CP(clk), .Q(\memory[6][40] ) );
  CFD1QXL \memory_reg[6][39]  ( .D(n1907), .CP(clk), .Q(\memory[6][39] ) );
  CFD1QXL \memory_reg[6][38]  ( .D(n1908), .CP(clk), .Q(\memory[6][38] ) );
  CFD1QXL \memory_reg[6][37]  ( .D(n1909), .CP(clk), .Q(\memory[6][37] ) );
  CFD1QXL \memory_reg[6][36]  ( .D(n1910), .CP(clk), .Q(\memory[6][36] ) );
  CFD1QXL \memory_reg[6][35]  ( .D(n1911), .CP(clk), .Q(\memory[6][35] ) );
  CFD1QXL \memory_reg[6][34]  ( .D(n1912), .CP(clk), .Q(\memory[6][34] ) );
  CFD1QXL \memory_reg[6][33]  ( .D(n1913), .CP(clk), .Q(\memory[6][33] ) );
  CFD1QXL \memory_reg[6][32]  ( .D(n1914), .CP(clk), .Q(\memory[6][32] ) );
  CFD1QXL \memory_reg[6][31]  ( .D(n1915), .CP(clk), .Q(\memory[6][31] ) );
  CFD1QXL \memory_reg[6][30]  ( .D(n1916), .CP(clk), .Q(\memory[6][30] ) );
  CFD1QXL \memory_reg[6][29]  ( .D(n1917), .CP(clk), .Q(\memory[6][29] ) );
  CFD1QXL \memory_reg[6][28]  ( .D(n1918), .CP(clk), .Q(\memory[6][28] ) );
  CFD1QXL \memory_reg[6][27]  ( .D(n1919), .CP(clk), .Q(\memory[6][27] ) );
  CFD1QXL \memory_reg[6][26]  ( .D(n1920), .CP(clk), .Q(\memory[6][26] ) );
  CFD1QXL \memory_reg[6][25]  ( .D(n1921), .CP(clk), .Q(\memory[6][25] ) );
  CFD1QXL \memory_reg[6][24]  ( .D(n1922), .CP(clk), .Q(\memory[6][24] ) );
  CFD1QXL \memory_reg[6][23]  ( .D(n1923), .CP(clk), .Q(\memory[6][23] ) );
  CFD1QXL \memory_reg[6][22]  ( .D(n1924), .CP(clk), .Q(\memory[6][22] ) );
  CFD1QXL \memory_reg[6][21]  ( .D(n1925), .CP(clk), .Q(\memory[6][21] ) );
  CFD1QXL \memory_reg[6][20]  ( .D(n1926), .CP(clk), .Q(\memory[6][20] ) );
  CFD1QXL \memory_reg[6][19]  ( .D(n1927), .CP(clk), .Q(\memory[6][19] ) );
  CFD1QXL \memory_reg[6][18]  ( .D(n1928), .CP(clk), .Q(\memory[6][18] ) );
  CFD1QXL \memory_reg[6][17]  ( .D(n1929), .CP(clk), .Q(\memory[6][17] ) );
  CFD1QXL \memory_reg[6][16]  ( .D(n1930), .CP(clk), .Q(\memory[6][16] ) );
  CFD1QXL \memory_reg[6][15]  ( .D(n1931), .CP(clk), .Q(\memory[6][15] ) );
  CFD1QXL \memory_reg[6][14]  ( .D(n1932), .CP(clk), .Q(\memory[6][14] ) );
  CFD1QXL \memory_reg[6][13]  ( .D(n1933), .CP(clk), .Q(\memory[6][13] ) );
  CFD1QXL \memory_reg[6][12]  ( .D(n1934), .CP(clk), .Q(\memory[6][12] ) );
  CFD1QXL \memory_reg[6][11]  ( .D(n1935), .CP(clk), .Q(\memory[6][11] ) );
  CFD1QXL \memory_reg[6][10]  ( .D(n1936), .CP(clk), .Q(\memory[6][10] ) );
  CFD1QXL \memory_reg[6][9]  ( .D(n1937), .CP(clk), .Q(\memory[6][9] ) );
  CFD1QXL \memory_reg[6][8]  ( .D(n1938), .CP(clk), .Q(\memory[6][8] ) );
  CFD1QXL \memory_reg[6][7]  ( .D(n1939), .CP(clk), .Q(\memory[6][7] ) );
  CFD1QXL \memory_reg[6][6]  ( .D(n1940), .CP(clk), .Q(\memory[6][6] ) );
  CFD1QXL \memory_reg[6][5]  ( .D(n1941), .CP(clk), .Q(\memory[6][5] ) );
  CFD1QXL \memory_reg[6][4]  ( .D(n1942), .CP(clk), .Q(\memory[6][4] ) );
  CFD1QXL \memory_reg[6][3]  ( .D(n1943), .CP(clk), .Q(\memory[6][3] ) );
  CFD1QXL \memory_reg[6][2]  ( .D(n1944), .CP(clk), .Q(\memory[6][2] ) );
  CFD1QXL \memory_reg[6][1]  ( .D(n1945), .CP(clk), .Q(\memory[6][1] ) );
  CFD1QXL \memory_reg[6][0]  ( .D(n1946), .CP(clk), .Q(\memory[6][0] ) );
  CFD1QXL \memory_reg[5][63]  ( .D(n1954), .CP(clk), .Q(\memory[5][63] ) );
  CFD1QXL \memory_reg[5][62]  ( .D(n1955), .CP(clk), .Q(\memory[5][62] ) );
  CFD1QXL \memory_reg[5][61]  ( .D(n1956), .CP(clk), .Q(\memory[5][61] ) );
  CFD1QXL \memory_reg[5][60]  ( .D(n1957), .CP(clk), .Q(\memory[5][60] ) );
  CFD1QXL \memory_reg[5][59]  ( .D(n1958), .CP(clk), .Q(\memory[5][59] ) );
  CFD1QXL \memory_reg[5][58]  ( .D(n1959), .CP(clk), .Q(\memory[5][58] ) );
  CFD1QXL \memory_reg[5][57]  ( .D(n1960), .CP(clk), .Q(\memory[5][57] ) );
  CFD1QXL \memory_reg[5][56]  ( .D(n1961), .CP(clk), .Q(\memory[5][56] ) );
  CFD1QXL \memory_reg[5][55]  ( .D(n1962), .CP(clk), .Q(\memory[5][55] ) );
  CFD1QXL \memory_reg[5][54]  ( .D(n1963), .CP(clk), .Q(\memory[5][54] ) );
  CFD1QXL \memory_reg[5][53]  ( .D(n1964), .CP(clk), .Q(\memory[5][53] ) );
  CFD1QXL \memory_reg[5][52]  ( .D(n1965), .CP(clk), .Q(\memory[5][52] ) );
  CFD1QXL \memory_reg[5][51]  ( .D(n1966), .CP(clk), .Q(\memory[5][51] ) );
  CFD1QXL \memory_reg[5][50]  ( .D(n1967), .CP(clk), .Q(\memory[5][50] ) );
  CFD1QXL \memory_reg[5][49]  ( .D(n1968), .CP(clk), .Q(\memory[5][49] ) );
  CFD1QXL \memory_reg[5][48]  ( .D(n1969), .CP(clk), .Q(\memory[5][48] ) );
  CFD1QXL \memory_reg[5][47]  ( .D(n1970), .CP(clk), .Q(\memory[5][47] ) );
  CFD1QXL \memory_reg[5][46]  ( .D(n1971), .CP(clk), .Q(\memory[5][46] ) );
  CFD1QXL \memory_reg[5][45]  ( .D(n1972), .CP(clk), .Q(\memory[5][45] ) );
  CFD1QXL \memory_reg[5][44]  ( .D(n1973), .CP(clk), .Q(\memory[5][44] ) );
  CFD1QXL \memory_reg[5][43]  ( .D(n1974), .CP(clk), .Q(\memory[5][43] ) );
  CFD1QXL \memory_reg[5][42]  ( .D(n1975), .CP(clk), .Q(\memory[5][42] ) );
  CFD1QXL \memory_reg[5][41]  ( .D(n1976), .CP(clk), .Q(\memory[5][41] ) );
  CFD1QXL \memory_reg[5][40]  ( .D(n1977), .CP(clk), .Q(\memory[5][40] ) );
  CFD1QXL \memory_reg[5][39]  ( .D(n1978), .CP(clk), .Q(\memory[5][39] ) );
  CFD1QXL \memory_reg[5][38]  ( .D(n1979), .CP(clk), .Q(\memory[5][38] ) );
  CFD1QXL \memory_reg[5][37]  ( .D(n1980), .CP(clk), .Q(\memory[5][37] ) );
  CFD1QXL \memory_reg[5][36]  ( .D(n1981), .CP(clk), .Q(\memory[5][36] ) );
  CFD1QXL \memory_reg[5][35]  ( .D(n1982), .CP(clk), .Q(\memory[5][35] ) );
  CFD1QXL \memory_reg[5][34]  ( .D(n1983), .CP(clk), .Q(\memory[5][34] ) );
  CFD1QXL \memory_reg[5][33]  ( .D(n1984), .CP(clk), .Q(\memory[5][33] ) );
  CFD1QXL \memory_reg[5][32]  ( .D(n1985), .CP(clk), .Q(\memory[5][32] ) );
  CFD1QXL \memory_reg[5][31]  ( .D(n1986), .CP(clk), .Q(\memory[5][31] ) );
  CFD1QXL \memory_reg[5][30]  ( .D(n1987), .CP(clk), .Q(\memory[5][30] ) );
  CFD1QXL \memory_reg[5][29]  ( .D(n1988), .CP(clk), .Q(\memory[5][29] ) );
  CFD1QXL \memory_reg[5][28]  ( .D(n1989), .CP(clk), .Q(\memory[5][28] ) );
  CFD1QXL \memory_reg[5][27]  ( .D(n1990), .CP(clk), .Q(\memory[5][27] ) );
  CFD1QXL \memory_reg[5][26]  ( .D(n1991), .CP(clk), .Q(\memory[5][26] ) );
  CFD1QXL \memory_reg[5][25]  ( .D(n1992), .CP(clk), .Q(\memory[5][25] ) );
  CFD1QXL \memory_reg[5][24]  ( .D(n1993), .CP(clk), .Q(\memory[5][24] ) );
  CFD1QXL \memory_reg[5][23]  ( .D(n1994), .CP(clk), .Q(\memory[5][23] ) );
  CFD1QXL \memory_reg[5][22]  ( .D(n1995), .CP(clk), .Q(\memory[5][22] ) );
  CFD1QXL \memory_reg[5][21]  ( .D(n1996), .CP(clk), .Q(\memory[5][21] ) );
  CFD1QXL \memory_reg[5][20]  ( .D(n1997), .CP(clk), .Q(\memory[5][20] ) );
  CFD1QXL \memory_reg[5][19]  ( .D(n1998), .CP(clk), .Q(\memory[5][19] ) );
  CFD1QXL \memory_reg[5][18]  ( .D(n1999), .CP(clk), .Q(\memory[5][18] ) );
  CFD1QXL \memory_reg[5][17]  ( .D(n2000), .CP(clk), .Q(\memory[5][17] ) );
  CFD1QXL \memory_reg[5][16]  ( .D(n2001), .CP(clk), .Q(\memory[5][16] ) );
  CFD1QXL \memory_reg[5][15]  ( .D(n2002), .CP(clk), .Q(\memory[5][15] ) );
  CFD1QXL \memory_reg[5][14]  ( .D(n2003), .CP(clk), .Q(\memory[5][14] ) );
  CFD1QXL \memory_reg[5][13]  ( .D(n2004), .CP(clk), .Q(\memory[5][13] ) );
  CFD1QXL \memory_reg[5][12]  ( .D(n2005), .CP(clk), .Q(\memory[5][12] ) );
  CFD1QXL \memory_reg[5][11]  ( .D(n2006), .CP(clk), .Q(\memory[5][11] ) );
  CFD1QXL \memory_reg[5][10]  ( .D(n2007), .CP(clk), .Q(\memory[5][10] ) );
  CFD1QXL \memory_reg[5][9]  ( .D(n2008), .CP(clk), .Q(\memory[5][9] ) );
  CFD1QXL \memory_reg[5][8]  ( .D(n2009), .CP(clk), .Q(\memory[5][8] ) );
  CFD1QXL \memory_reg[5][7]  ( .D(n2010), .CP(clk), .Q(\memory[5][7] ) );
  CFD1QXL \memory_reg[5][6]  ( .D(n2011), .CP(clk), .Q(\memory[5][6] ) );
  CFD1QXL \memory_reg[5][5]  ( .D(n2012), .CP(clk), .Q(\memory[5][5] ) );
  CFD1QXL \memory_reg[5][4]  ( .D(n2013), .CP(clk), .Q(\memory[5][4] ) );
  CFD1QXL \memory_reg[5][3]  ( .D(n2014), .CP(clk), .Q(\memory[5][3] ) );
  CFD1QXL \memory_reg[5][2]  ( .D(n2015), .CP(clk), .Q(\memory[5][2] ) );
  CFD1QXL \memory_reg[5][1]  ( .D(n2016), .CP(clk), .Q(\memory[5][1] ) );
  CFD1QXL \memory_reg[5][0]  ( .D(n2017), .CP(clk), .Q(\memory[5][0] ) );
  CFD1QXL \memory_reg[4][63]  ( .D(n2025), .CP(clk), .Q(\memory[4][63] ) );
  CFD1QXL \memory_reg[4][62]  ( .D(n2026), .CP(clk), .Q(\memory[4][62] ) );
  CFD1QXL \memory_reg[4][61]  ( .D(n2027), .CP(clk), .Q(\memory[4][61] ) );
  CFD1QXL \memory_reg[4][60]  ( .D(n2028), .CP(clk), .Q(\memory[4][60] ) );
  CFD1QXL \memory_reg[4][59]  ( .D(n2029), .CP(clk), .Q(\memory[4][59] ) );
  CFD1QXL \memory_reg[4][58]  ( .D(n2030), .CP(clk), .Q(\memory[4][58] ) );
  CFD1QXL \memory_reg[4][57]  ( .D(n2031), .CP(clk), .Q(\memory[4][57] ) );
  CFD1QXL \memory_reg[4][56]  ( .D(n2032), .CP(clk), .Q(\memory[4][56] ) );
  CFD1QXL \memory_reg[4][55]  ( .D(n2033), .CP(clk), .Q(\memory[4][55] ) );
  CFD1QXL \memory_reg[4][54]  ( .D(n2034), .CP(clk), .Q(\memory[4][54] ) );
  CFD1QXL \memory_reg[4][53]  ( .D(n2035), .CP(clk), .Q(\memory[4][53] ) );
  CFD1QXL \memory_reg[4][52]  ( .D(n2036), .CP(clk), .Q(\memory[4][52] ) );
  CFD1QXL \memory_reg[4][51]  ( .D(n2037), .CP(clk), .Q(\memory[4][51] ) );
  CFD1QXL \memory_reg[4][50]  ( .D(n2038), .CP(clk), .Q(\memory[4][50] ) );
  CFD1QXL \memory_reg[4][49]  ( .D(n2039), .CP(clk), .Q(\memory[4][49] ) );
  CFD1QXL \memory_reg[4][48]  ( .D(n2040), .CP(clk), .Q(\memory[4][48] ) );
  CFD1QXL \memory_reg[4][47]  ( .D(n2041), .CP(clk), .Q(\memory[4][47] ) );
  CFD1QXL \memory_reg[4][46]  ( .D(n2042), .CP(clk), .Q(\memory[4][46] ) );
  CFD1QXL \memory_reg[4][45]  ( .D(n2043), .CP(clk), .Q(\memory[4][45] ) );
  CFD1QXL \memory_reg[4][44]  ( .D(n2044), .CP(clk), .Q(\memory[4][44] ) );
  CFD1QXL \memory_reg[4][43]  ( .D(n2045), .CP(clk), .Q(\memory[4][43] ) );
  CFD1QXL \memory_reg[4][42]  ( .D(n2046), .CP(clk), .Q(\memory[4][42] ) );
  CFD1QXL \memory_reg[4][41]  ( .D(n2047), .CP(clk), .Q(\memory[4][41] ) );
  CFD1QXL \memory_reg[4][40]  ( .D(n2048), .CP(clk), .Q(\memory[4][40] ) );
  CFD1QXL \memory_reg[4][39]  ( .D(n2049), .CP(clk), .Q(\memory[4][39] ) );
  CFD1QXL \memory_reg[4][38]  ( .D(n2050), .CP(clk), .Q(\memory[4][38] ) );
  CFD1QXL \memory_reg[4][37]  ( .D(n2051), .CP(clk), .Q(\memory[4][37] ) );
  CFD1QXL \memory_reg[4][36]  ( .D(n2052), .CP(clk), .Q(\memory[4][36] ) );
  CFD1QXL \memory_reg[4][35]  ( .D(n2053), .CP(clk), .Q(\memory[4][35] ) );
  CFD1QXL \memory_reg[4][34]  ( .D(n2054), .CP(clk), .Q(\memory[4][34] ) );
  CFD1QXL \memory_reg[4][33]  ( .D(n2055), .CP(clk), .Q(\memory[4][33] ) );
  CFD1QXL \memory_reg[4][32]  ( .D(n2056), .CP(clk), .Q(\memory[4][32] ) );
  CFD1QXL \memory_reg[4][31]  ( .D(n2057), .CP(clk), .Q(\memory[4][31] ) );
  CFD1QXL \memory_reg[4][30]  ( .D(n2058), .CP(clk), .Q(\memory[4][30] ) );
  CFD1QXL \memory_reg[4][29]  ( .D(n2059), .CP(clk), .Q(\memory[4][29] ) );
  CFD1QXL \memory_reg[4][28]  ( .D(n2060), .CP(clk), .Q(\memory[4][28] ) );
  CFD1QXL \memory_reg[4][27]  ( .D(n2061), .CP(clk), .Q(\memory[4][27] ) );
  CFD1QXL \memory_reg[4][26]  ( .D(n2062), .CP(clk), .Q(\memory[4][26] ) );
  CFD1QXL \memory_reg[4][25]  ( .D(n2063), .CP(clk), .Q(\memory[4][25] ) );
  CFD1QXL \memory_reg[4][24]  ( .D(n2064), .CP(clk), .Q(\memory[4][24] ) );
  CFD1QXL \memory_reg[4][23]  ( .D(n2065), .CP(clk), .Q(\memory[4][23] ) );
  CFD1QXL \memory_reg[4][22]  ( .D(n2066), .CP(clk), .Q(\memory[4][22] ) );
  CFD1QXL \memory_reg[4][21]  ( .D(n2067), .CP(clk), .Q(\memory[4][21] ) );
  CFD1QXL \memory_reg[4][20]  ( .D(n2068), .CP(clk), .Q(\memory[4][20] ) );
  CFD1QXL \memory_reg[4][19]  ( .D(n2069), .CP(clk), .Q(\memory[4][19] ) );
  CFD1QXL \memory_reg[4][18]  ( .D(n2070), .CP(clk), .Q(\memory[4][18] ) );
  CFD1QXL \memory_reg[4][17]  ( .D(n2071), .CP(clk), .Q(\memory[4][17] ) );
  CFD1QXL \memory_reg[4][16]  ( .D(n2072), .CP(clk), .Q(\memory[4][16] ) );
  CFD1QXL \memory_reg[4][15]  ( .D(n2073), .CP(clk), .Q(\memory[4][15] ) );
  CFD1QXL \memory_reg[4][14]  ( .D(n2074), .CP(clk), .Q(\memory[4][14] ) );
  CFD1QXL \memory_reg[4][13]  ( .D(n2075), .CP(clk), .Q(\memory[4][13] ) );
  CFD1QXL \memory_reg[4][12]  ( .D(n2076), .CP(clk), .Q(\memory[4][12] ) );
  CFD1QXL \memory_reg[4][11]  ( .D(n2077), .CP(clk), .Q(\memory[4][11] ) );
  CFD1QXL \memory_reg[4][10]  ( .D(n2078), .CP(clk), .Q(\memory[4][10] ) );
  CFD1QXL \memory_reg[4][9]  ( .D(n2079), .CP(clk), .Q(\memory[4][9] ) );
  CFD1QXL \memory_reg[4][8]  ( .D(n2080), .CP(clk), .Q(\memory[4][8] ) );
  CFD1QXL \memory_reg[4][7]  ( .D(n2081), .CP(clk), .Q(\memory[4][7] ) );
  CFD1QXL \memory_reg[4][6]  ( .D(n2082), .CP(clk), .Q(\memory[4][6] ) );
  CFD1QXL \memory_reg[4][5]  ( .D(n2083), .CP(clk), .Q(\memory[4][5] ) );
  CFD1QXL \memory_reg[4][4]  ( .D(n2084), .CP(clk), .Q(\memory[4][4] ) );
  CFD1QXL \memory_reg[4][3]  ( .D(n2085), .CP(clk), .Q(\memory[4][3] ) );
  CFD1QXL \memory_reg[4][2]  ( .D(n2086), .CP(clk), .Q(\memory[4][2] ) );
  CFD1QXL \memory_reg[4][1]  ( .D(n2087), .CP(clk), .Q(\memory[4][1] ) );
  CFD1QXL \memory_reg[4][0]  ( .D(n2088), .CP(clk), .Q(\memory[4][0] ) );
  CFD1QXL \memory_reg[3][63]  ( .D(n2096), .CP(clk), .Q(\memory[3][63] ) );
  CFD1QXL \memory_reg[3][62]  ( .D(n2097), .CP(clk), .Q(\memory[3][62] ) );
  CFD1QXL \memory_reg[3][61]  ( .D(n2098), .CP(clk), .Q(\memory[3][61] ) );
  CFD1QXL \memory_reg[3][60]  ( .D(n2099), .CP(clk), .Q(\memory[3][60] ) );
  CFD1QXL \memory_reg[3][59]  ( .D(n2100), .CP(clk), .Q(\memory[3][59] ) );
  CFD1QXL \memory_reg[3][58]  ( .D(n2101), .CP(clk), .Q(\memory[3][58] ) );
  CFD1QXL \memory_reg[3][57]  ( .D(n2102), .CP(clk), .Q(\memory[3][57] ) );
  CFD1QXL \memory_reg[3][56]  ( .D(n2103), .CP(clk), .Q(\memory[3][56] ) );
  CFD1QXL \memory_reg[3][55]  ( .D(n2104), .CP(clk), .Q(\memory[3][55] ) );
  CFD1QXL \memory_reg[3][54]  ( .D(n2105), .CP(clk), .Q(\memory[3][54] ) );
  CFD1QXL \memory_reg[3][53]  ( .D(n2106), .CP(clk), .Q(\memory[3][53] ) );
  CFD1QXL \memory_reg[3][52]  ( .D(n2107), .CP(clk), .Q(\memory[3][52] ) );
  CFD1QXL \memory_reg[3][51]  ( .D(n2108), .CP(clk), .Q(\memory[3][51] ) );
  CFD1QXL \memory_reg[3][50]  ( .D(n2109), .CP(clk), .Q(\memory[3][50] ) );
  CFD1QXL \memory_reg[3][49]  ( .D(n2110), .CP(clk), .Q(\memory[3][49] ) );
  CFD1QXL \memory_reg[3][48]  ( .D(n2111), .CP(clk), .Q(\memory[3][48] ) );
  CFD1QXL \memory_reg[3][47]  ( .D(n2112), .CP(clk), .Q(\memory[3][47] ) );
  CFD1QXL \memory_reg[3][46]  ( .D(n2113), .CP(clk), .Q(\memory[3][46] ) );
  CFD1QXL \memory_reg[3][45]  ( .D(n2114), .CP(clk), .Q(\memory[3][45] ) );
  CFD1QXL \memory_reg[3][44]  ( .D(n2115), .CP(clk), .Q(\memory[3][44] ) );
  CFD1QXL \memory_reg[3][43]  ( .D(n2116), .CP(clk), .Q(\memory[3][43] ) );
  CFD1QXL \memory_reg[3][42]  ( .D(n2117), .CP(clk), .Q(\memory[3][42] ) );
  CFD1QXL \memory_reg[3][41]  ( .D(n2118), .CP(clk), .Q(\memory[3][41] ) );
  CFD1QXL \memory_reg[3][40]  ( .D(n2119), .CP(clk), .Q(\memory[3][40] ) );
  CFD1QXL \memory_reg[3][39]  ( .D(n2120), .CP(clk), .Q(\memory[3][39] ) );
  CFD1QXL \memory_reg[3][38]  ( .D(n2121), .CP(clk), .Q(\memory[3][38] ) );
  CFD1QXL \memory_reg[3][37]  ( .D(n2122), .CP(clk), .Q(\memory[3][37] ) );
  CFD1QXL \memory_reg[3][36]  ( .D(n2123), .CP(clk), .Q(\memory[3][36] ) );
  CFD1QXL \memory_reg[3][35]  ( .D(n2124), .CP(clk), .Q(\memory[3][35] ) );
  CFD1QXL \memory_reg[3][34]  ( .D(n2125), .CP(clk), .Q(\memory[3][34] ) );
  CFD1QXL \memory_reg[3][33]  ( .D(n2126), .CP(clk), .Q(\memory[3][33] ) );
  CFD1QXL \memory_reg[3][32]  ( .D(n2127), .CP(clk), .Q(\memory[3][32] ) );
  CFD1QXL \memory_reg[3][31]  ( .D(n2128), .CP(clk), .Q(\memory[3][31] ) );
  CFD1QXL \memory_reg[3][30]  ( .D(n2129), .CP(clk), .Q(\memory[3][30] ) );
  CFD1QXL \memory_reg[3][29]  ( .D(n2130), .CP(clk), .Q(\memory[3][29] ) );
  CFD1QXL \memory_reg[3][28]  ( .D(n2131), .CP(clk), .Q(\memory[3][28] ) );
  CFD1QXL \memory_reg[3][27]  ( .D(n2132), .CP(clk), .Q(\memory[3][27] ) );
  CFD1QXL \memory_reg[3][26]  ( .D(n2133), .CP(clk), .Q(\memory[3][26] ) );
  CFD1QXL \memory_reg[3][25]  ( .D(n2134), .CP(clk), .Q(\memory[3][25] ) );
  CFD1QXL \memory_reg[3][24]  ( .D(n2135), .CP(clk), .Q(\memory[3][24] ) );
  CFD1QXL \memory_reg[3][23]  ( .D(n2136), .CP(clk), .Q(\memory[3][23] ) );
  CFD1QXL \memory_reg[3][22]  ( .D(n2137), .CP(clk), .Q(\memory[3][22] ) );
  CFD1QXL \memory_reg[3][21]  ( .D(n2138), .CP(clk), .Q(\memory[3][21] ) );
  CFD1QXL \memory_reg[3][20]  ( .D(n2139), .CP(clk), .Q(\memory[3][20] ) );
  CFD1QXL \memory_reg[3][19]  ( .D(n2140), .CP(clk), .Q(\memory[3][19] ) );
  CFD1QXL \memory_reg[3][18]  ( .D(n2141), .CP(clk), .Q(\memory[3][18] ) );
  CFD1QXL \memory_reg[3][17]  ( .D(n2142), .CP(clk), .Q(\memory[3][17] ) );
  CFD1QXL \memory_reg[3][16]  ( .D(n2143), .CP(clk), .Q(\memory[3][16] ) );
  CFD1QXL \memory_reg[3][15]  ( .D(n2144), .CP(clk), .Q(\memory[3][15] ) );
  CFD1QXL \memory_reg[3][14]  ( .D(n2145), .CP(clk), .Q(\memory[3][14] ) );
  CFD1QXL \memory_reg[3][13]  ( .D(n2146), .CP(clk), .Q(\memory[3][13] ) );
  CFD1QXL \memory_reg[3][12]  ( .D(n2147), .CP(clk), .Q(\memory[3][12] ) );
  CFD1QXL \memory_reg[3][11]  ( .D(n2148), .CP(clk), .Q(\memory[3][11] ) );
  CFD1QXL \memory_reg[3][10]  ( .D(n2149), .CP(clk), .Q(\memory[3][10] ) );
  CFD1QXL \memory_reg[3][9]  ( .D(n2150), .CP(clk), .Q(\memory[3][9] ) );
  CFD1QXL \memory_reg[3][8]  ( .D(n2151), .CP(clk), .Q(\memory[3][8] ) );
  CFD1QXL \memory_reg[3][7]  ( .D(n2152), .CP(clk), .Q(\memory[3][7] ) );
  CFD1QXL \memory_reg[3][6]  ( .D(n2153), .CP(clk), .Q(\memory[3][6] ) );
  CFD1QXL \memory_reg[3][5]  ( .D(n2154), .CP(clk), .Q(\memory[3][5] ) );
  CFD1QXL \memory_reg[3][4]  ( .D(n2155), .CP(clk), .Q(\memory[3][4] ) );
  CFD1QXL \memory_reg[3][3]  ( .D(n2156), .CP(clk), .Q(\memory[3][3] ) );
  CFD1QXL \memory_reg[3][2]  ( .D(n2157), .CP(clk), .Q(\memory[3][2] ) );
  CFD1QXL \memory_reg[3][1]  ( .D(n2158), .CP(clk), .Q(\memory[3][1] ) );
  CFD1QXL \memory_reg[3][0]  ( .D(n2159), .CP(clk), .Q(\memory[3][0] ) );
  CFD1QXL \memory_reg[2][63]  ( .D(n2167), .CP(clk), .Q(\memory[2][63] ) );
  CFD1QXL \memory_reg[2][62]  ( .D(n2168), .CP(clk), .Q(\memory[2][62] ) );
  CFD1QXL \memory_reg[2][61]  ( .D(n2169), .CP(clk), .Q(\memory[2][61] ) );
  CFD1QXL \memory_reg[2][60]  ( .D(n2170), .CP(clk), .Q(\memory[2][60] ) );
  CFD1QXL \memory_reg[2][59]  ( .D(n2171), .CP(clk), .Q(\memory[2][59] ) );
  CFD1QXL \memory_reg[2][58]  ( .D(n2172), .CP(clk), .Q(\memory[2][58] ) );
  CFD1QXL \memory_reg[2][57]  ( .D(n2173), .CP(clk), .Q(\memory[2][57] ) );
  CFD1QXL \memory_reg[2][56]  ( .D(n2174), .CP(clk), .Q(\memory[2][56] ) );
  CFD1QXL \memory_reg[2][55]  ( .D(n2175), .CP(clk), .Q(\memory[2][55] ) );
  CFD1QXL \memory_reg[2][54]  ( .D(n2176), .CP(clk), .Q(\memory[2][54] ) );
  CFD1QXL \memory_reg[2][53]  ( .D(n2177), .CP(clk), .Q(\memory[2][53] ) );
  CFD1QXL \memory_reg[2][52]  ( .D(n2178), .CP(clk), .Q(\memory[2][52] ) );
  CFD1QXL \memory_reg[2][51]  ( .D(n2179), .CP(clk), .Q(\memory[2][51] ) );
  CFD1QXL \memory_reg[2][50]  ( .D(n2180), .CP(clk), .Q(\memory[2][50] ) );
  CFD1QXL \memory_reg[2][49]  ( .D(n2181), .CP(clk), .Q(\memory[2][49] ) );
  CFD1QXL \memory_reg[2][48]  ( .D(n2182), .CP(clk), .Q(\memory[2][48] ) );
  CFD1QXL \memory_reg[2][47]  ( .D(n2183), .CP(clk), .Q(\memory[2][47] ) );
  CFD1QXL \memory_reg[2][46]  ( .D(n2184), .CP(clk), .Q(\memory[2][46] ) );
  CFD1QXL \memory_reg[2][45]  ( .D(n2185), .CP(clk), .Q(\memory[2][45] ) );
  CFD1QXL \memory_reg[2][44]  ( .D(n2186), .CP(clk), .Q(\memory[2][44] ) );
  CFD1QXL \memory_reg[2][43]  ( .D(n2187), .CP(clk), .Q(\memory[2][43] ) );
  CFD1QXL \memory_reg[2][42]  ( .D(n2188), .CP(clk), .Q(\memory[2][42] ) );
  CFD1QXL \memory_reg[2][41]  ( .D(n2189), .CP(clk), .Q(\memory[2][41] ) );
  CFD1QXL \memory_reg[2][40]  ( .D(n2190), .CP(clk), .Q(\memory[2][40] ) );
  CFD1QXL \memory_reg[2][39]  ( .D(n2191), .CP(clk), .Q(\memory[2][39] ) );
  CFD1QXL \memory_reg[2][38]  ( .D(n2192), .CP(clk), .Q(\memory[2][38] ) );
  CFD1QXL \memory_reg[2][37]  ( .D(n2193), .CP(clk), .Q(\memory[2][37] ) );
  CFD1QXL \memory_reg[2][36]  ( .D(n2194), .CP(clk), .Q(\memory[2][36] ) );
  CFD1QXL \memory_reg[2][35]  ( .D(n2195), .CP(clk), .Q(\memory[2][35] ) );
  CFD1QXL \memory_reg[2][34]  ( .D(n2196), .CP(clk), .Q(\memory[2][34] ) );
  CFD1QXL \memory_reg[2][33]  ( .D(n2197), .CP(clk), .Q(\memory[2][33] ) );
  CFD1QXL \memory_reg[2][32]  ( .D(n2198), .CP(clk), .Q(\memory[2][32] ) );
  CFD1QXL \memory_reg[2][31]  ( .D(n2199), .CP(clk), .Q(\memory[2][31] ) );
  CFD1QXL \memory_reg[2][30]  ( .D(n2200), .CP(clk), .Q(\memory[2][30] ) );
  CFD1QXL \memory_reg[2][29]  ( .D(n2201), .CP(clk), .Q(\memory[2][29] ) );
  CFD1QXL \memory_reg[2][28]  ( .D(n2202), .CP(clk), .Q(\memory[2][28] ) );
  CFD1QXL \memory_reg[2][27]  ( .D(n2203), .CP(clk), .Q(\memory[2][27] ) );
  CFD1QXL \memory_reg[2][26]  ( .D(n2204), .CP(clk), .Q(\memory[2][26] ) );
  CFD1QXL \memory_reg[2][25]  ( .D(n2205), .CP(clk), .Q(\memory[2][25] ) );
  CFD1QXL \memory_reg[2][24]  ( .D(n2206), .CP(clk), .Q(\memory[2][24] ) );
  CFD1QXL \memory_reg[2][23]  ( .D(n2207), .CP(clk), .Q(\memory[2][23] ) );
  CFD1QXL \memory_reg[2][22]  ( .D(n2208), .CP(clk), .Q(\memory[2][22] ) );
  CFD1QXL \memory_reg[2][21]  ( .D(n2209), .CP(clk), .Q(\memory[2][21] ) );
  CFD1QXL \memory_reg[2][20]  ( .D(n2210), .CP(clk), .Q(\memory[2][20] ) );
  CFD1QXL \memory_reg[2][19]  ( .D(n2211), .CP(clk), .Q(\memory[2][19] ) );
  CFD1QXL \memory_reg[2][18]  ( .D(n2212), .CP(clk), .Q(\memory[2][18] ) );
  CFD1QXL \memory_reg[2][17]  ( .D(n2213), .CP(clk), .Q(\memory[2][17] ) );
  CFD1QXL \memory_reg[2][16]  ( .D(n2214), .CP(clk), .Q(\memory[2][16] ) );
  CFD1QXL \memory_reg[2][15]  ( .D(n2215), .CP(clk), .Q(\memory[2][15] ) );
  CFD1QXL \memory_reg[2][14]  ( .D(n2216), .CP(clk), .Q(\memory[2][14] ) );
  CFD1QXL \memory_reg[2][13]  ( .D(n2217), .CP(clk), .Q(\memory[2][13] ) );
  CFD1QXL \memory_reg[2][12]  ( .D(n2218), .CP(clk), .Q(\memory[2][12] ) );
  CFD1QXL \memory_reg[2][11]  ( .D(n2219), .CP(clk), .Q(\memory[2][11] ) );
  CFD1QXL \memory_reg[2][10]  ( .D(n2220), .CP(clk), .Q(\memory[2][10] ) );
  CFD1QXL \memory_reg[2][9]  ( .D(n2221), .CP(clk), .Q(\memory[2][9] ) );
  CFD1QXL \memory_reg[2][8]  ( .D(n2222), .CP(clk), .Q(\memory[2][8] ) );
  CFD1QXL \memory_reg[2][7]  ( .D(n2223), .CP(clk), .Q(\memory[2][7] ) );
  CFD1QXL \memory_reg[2][6]  ( .D(n2224), .CP(clk), .Q(\memory[2][6] ) );
  CFD1QXL \memory_reg[2][5]  ( .D(n2225), .CP(clk), .Q(\memory[2][5] ) );
  CFD1QXL \memory_reg[2][4]  ( .D(n2226), .CP(clk), .Q(\memory[2][4] ) );
  CFD1QXL \memory_reg[2][3]  ( .D(n2227), .CP(clk), .Q(\memory[2][3] ) );
  CFD1QXL \memory_reg[2][2]  ( .D(n2228), .CP(clk), .Q(\memory[2][2] ) );
  CFD1QXL \memory_reg[2][1]  ( .D(n2229), .CP(clk), .Q(\memory[2][1] ) );
  CFD1QXL \memory_reg[2][0]  ( .D(n2230), .CP(clk), .Q(\memory[2][0] ) );
  CFD1QXL \memory_reg[1][63]  ( .D(n2238), .CP(clk), .Q(\memory[1][63] ) );
  CFD1QXL \memory_reg[1][62]  ( .D(n2239), .CP(clk), .Q(\memory[1][62] ) );
  CFD1QXL \memory_reg[1][61]  ( .D(n2240), .CP(clk), .Q(\memory[1][61] ) );
  CFD1QXL \memory_reg[1][60]  ( .D(n2241), .CP(clk), .Q(\memory[1][60] ) );
  CFD1QXL \memory_reg[1][59]  ( .D(n2242), .CP(clk), .Q(\memory[1][59] ) );
  CFD1QXL \memory_reg[1][58]  ( .D(n2243), .CP(clk), .Q(\memory[1][58] ) );
  CFD1QXL \memory_reg[1][57]  ( .D(n2244), .CP(clk), .Q(\memory[1][57] ) );
  CFD1QXL \memory_reg[1][56]  ( .D(n2245), .CP(clk), .Q(\memory[1][56] ) );
  CFD1QXL \memory_reg[1][55]  ( .D(n2246), .CP(clk), .Q(\memory[1][55] ) );
  CFD1QXL \memory_reg[1][54]  ( .D(n2247), .CP(clk), .Q(\memory[1][54] ) );
  CFD1QXL \memory_reg[1][53]  ( .D(n2248), .CP(clk), .Q(\memory[1][53] ) );
  CFD1QXL \memory_reg[1][52]  ( .D(n2249), .CP(clk), .Q(\memory[1][52] ) );
  CFD1QXL \memory_reg[1][51]  ( .D(n2250), .CP(clk), .Q(\memory[1][51] ) );
  CFD1QXL \memory_reg[1][50]  ( .D(n2251), .CP(clk), .Q(\memory[1][50] ) );
  CFD1QXL \memory_reg[1][49]  ( .D(n2252), .CP(clk), .Q(\memory[1][49] ) );
  CFD1QXL \memory_reg[1][48]  ( .D(n2253), .CP(clk), .Q(\memory[1][48] ) );
  CFD1QXL \memory_reg[1][47]  ( .D(n2254), .CP(clk), .Q(\memory[1][47] ) );
  CFD1QXL \memory_reg[1][46]  ( .D(n2255), .CP(clk), .Q(\memory[1][46] ) );
  CFD1QXL \memory_reg[1][45]  ( .D(n2256), .CP(clk), .Q(\memory[1][45] ) );
  CFD1QXL \memory_reg[1][44]  ( .D(n2257), .CP(clk), .Q(\memory[1][44] ) );
  CFD1QXL \memory_reg[1][43]  ( .D(n2258), .CP(clk), .Q(\memory[1][43] ) );
  CFD1QXL \memory_reg[1][42]  ( .D(n2259), .CP(clk), .Q(\memory[1][42] ) );
  CFD1QXL \memory_reg[1][41]  ( .D(n2260), .CP(clk), .Q(\memory[1][41] ) );
  CFD1QXL \memory_reg[1][40]  ( .D(n2261), .CP(clk), .Q(\memory[1][40] ) );
  CFD1QXL \memory_reg[1][39]  ( .D(n2262), .CP(clk), .Q(\memory[1][39] ) );
  CFD1QXL \memory_reg[1][38]  ( .D(n2263), .CP(clk), .Q(\memory[1][38] ) );
  CFD1QXL \memory_reg[1][37]  ( .D(n2264), .CP(clk), .Q(\memory[1][37] ) );
  CFD1QXL \memory_reg[1][36]  ( .D(n2265), .CP(clk), .Q(\memory[1][36] ) );
  CFD1QXL \memory_reg[1][35]  ( .D(n2266), .CP(clk), .Q(\memory[1][35] ) );
  CFD1QXL \memory_reg[1][34]  ( .D(n2267), .CP(clk), .Q(\memory[1][34] ) );
  CFD1QXL \memory_reg[1][33]  ( .D(n2268), .CP(clk), .Q(\memory[1][33] ) );
  CFD1QXL \memory_reg[1][32]  ( .D(n2269), .CP(clk), .Q(\memory[1][32] ) );
  CFD1QXL \memory_reg[1][31]  ( .D(n2270), .CP(clk), .Q(\memory[1][31] ) );
  CFD1QXL \memory_reg[1][30]  ( .D(n2271), .CP(clk), .Q(\memory[1][30] ) );
  CFD1QXL \memory_reg[1][29]  ( .D(n2272), .CP(clk), .Q(\memory[1][29] ) );
  CFD1QXL \memory_reg[1][28]  ( .D(n2273), .CP(clk), .Q(\memory[1][28] ) );
  CFD1QXL \memory_reg[1][27]  ( .D(n2274), .CP(clk), .Q(\memory[1][27] ) );
  CFD1QXL \memory_reg[1][26]  ( .D(n2275), .CP(clk), .Q(\memory[1][26] ) );
  CFD1QXL \memory_reg[1][25]  ( .D(n2276), .CP(clk), .Q(\memory[1][25] ) );
  CFD1QXL \memory_reg[1][24]  ( .D(n2277), .CP(clk), .Q(\memory[1][24] ) );
  CFD1QXL \memory_reg[1][23]  ( .D(n2278), .CP(clk), .Q(\memory[1][23] ) );
  CFD1QXL \memory_reg[1][22]  ( .D(n2279), .CP(clk), .Q(\memory[1][22] ) );
  CFD1QXL \memory_reg[1][21]  ( .D(n2280), .CP(clk), .Q(\memory[1][21] ) );
  CFD1QXL \memory_reg[1][20]  ( .D(n2281), .CP(clk), .Q(\memory[1][20] ) );
  CFD1QXL \memory_reg[1][19]  ( .D(n2282), .CP(clk), .Q(\memory[1][19] ) );
  CFD1QXL \memory_reg[1][18]  ( .D(n2283), .CP(clk), .Q(\memory[1][18] ) );
  CFD1QXL \memory_reg[1][17]  ( .D(n2284), .CP(clk), .Q(\memory[1][17] ) );
  CFD1QXL \memory_reg[1][16]  ( .D(n2285), .CP(clk), .Q(\memory[1][16] ) );
  CFD1QXL \memory_reg[1][15]  ( .D(n2286), .CP(clk), .Q(\memory[1][15] ) );
  CFD1QXL \memory_reg[1][14]  ( .D(n2287), .CP(clk), .Q(\memory[1][14] ) );
  CFD1QXL \memory_reg[1][13]  ( .D(n2288), .CP(clk), .Q(\memory[1][13] ) );
  CFD1QXL \memory_reg[1][12]  ( .D(n2289), .CP(clk), .Q(\memory[1][12] ) );
  CFD1QXL \memory_reg[1][11]  ( .D(n2290), .CP(clk), .Q(\memory[1][11] ) );
  CFD1QXL \memory_reg[1][10]  ( .D(n2291), .CP(clk), .Q(\memory[1][10] ) );
  CFD1QXL \memory_reg[1][9]  ( .D(n2292), .CP(clk), .Q(\memory[1][9] ) );
  CFD1QXL \memory_reg[1][8]  ( .D(n2293), .CP(clk), .Q(\memory[1][8] ) );
  CFD1QXL \memory_reg[1][7]  ( .D(n2294), .CP(clk), .Q(\memory[1][7] ) );
  CFD1QXL \memory_reg[1][6]  ( .D(n2295), .CP(clk), .Q(\memory[1][6] ) );
  CFD1QXL \memory_reg[1][5]  ( .D(n2296), .CP(clk), .Q(\memory[1][5] ) );
  CFD1QXL \memory_reg[1][4]  ( .D(n2297), .CP(clk), .Q(\memory[1][4] ) );
  CFD1QXL \memory_reg[1][3]  ( .D(n2298), .CP(clk), .Q(\memory[1][3] ) );
  CFD1QXL \memory_reg[1][2]  ( .D(n2299), .CP(clk), .Q(\memory[1][2] ) );
  CFD1QXL \memory_reg[1][1]  ( .D(n2300), .CP(clk), .Q(\memory[1][1] ) );
  CFD1QXL \memory_reg[1][0]  ( .D(n2301), .CP(clk), .Q(\memory[1][0] ) );
  CFD1QXL \memory_reg[0][63]  ( .D(n2309), .CP(clk), .Q(\memory[0][63] ) );
  CFD1QXL \memory_reg[0][62]  ( .D(n2310), .CP(clk), .Q(\memory[0][62] ) );
  CFD1QXL \memory_reg[0][61]  ( .D(n2311), .CP(clk), .Q(\memory[0][61] ) );
  CFD1QXL \memory_reg[0][60]  ( .D(n2312), .CP(clk), .Q(\memory[0][60] ) );
  CFD1QXL \memory_reg[0][59]  ( .D(n2313), .CP(clk), .Q(\memory[0][59] ) );
  CFD1QXL \memory_reg[0][58]  ( .D(n2314), .CP(clk), .Q(\memory[0][58] ) );
  CFD1QXL \memory_reg[0][57]  ( .D(n2315), .CP(clk), .Q(\memory[0][57] ) );
  CFD1QXL \memory_reg[0][56]  ( .D(n2316), .CP(clk), .Q(\memory[0][56] ) );
  CFD1QXL \memory_reg[0][55]  ( .D(n2317), .CP(clk), .Q(\memory[0][55] ) );
  CFD1QXL \memory_reg[0][54]  ( .D(n2318), .CP(clk), .Q(\memory[0][54] ) );
  CFD1QXL \memory_reg[0][53]  ( .D(n2319), .CP(clk), .Q(\memory[0][53] ) );
  CFD1QXL \memory_reg[0][52]  ( .D(n2320), .CP(clk), .Q(\memory[0][52] ) );
  CFD1QXL \memory_reg[0][51]  ( .D(n2321), .CP(clk), .Q(\memory[0][51] ) );
  CFD1QXL \memory_reg[0][50]  ( .D(n2322), .CP(clk), .Q(\memory[0][50] ) );
  CFD1QXL \memory_reg[0][49]  ( .D(n2323), .CP(clk), .Q(\memory[0][49] ) );
  CFD1QXL \memory_reg[0][48]  ( .D(n2324), .CP(clk), .Q(\memory[0][48] ) );
  CFD1QXL \memory_reg[0][47]  ( .D(n2325), .CP(clk), .Q(\memory[0][47] ) );
  CFD1QXL \memory_reg[0][46]  ( .D(n2326), .CP(clk), .Q(\memory[0][46] ) );
  CFD1QXL \memory_reg[0][45]  ( .D(n2327), .CP(clk), .Q(\memory[0][45] ) );
  CFD1QXL \memory_reg[0][44]  ( .D(n2328), .CP(clk), .Q(\memory[0][44] ) );
  CFD1QXL \memory_reg[0][43]  ( .D(n2329), .CP(clk), .Q(\memory[0][43] ) );
  CFD1QXL \memory_reg[0][42]  ( .D(n2330), .CP(clk), .Q(\memory[0][42] ) );
  CFD1QXL \memory_reg[0][41]  ( .D(n2331), .CP(clk), .Q(\memory[0][41] ) );
  CFD1QXL \memory_reg[0][40]  ( .D(n2332), .CP(clk), .Q(\memory[0][40] ) );
  CFD1QXL \memory_reg[0][39]  ( .D(n2333), .CP(clk), .Q(\memory[0][39] ) );
  CFD1QXL \memory_reg[0][38]  ( .D(n2334), .CP(clk), .Q(\memory[0][38] ) );
  CFD1QXL \memory_reg[0][37]  ( .D(n2335), .CP(clk), .Q(\memory[0][37] ) );
  CFD1QXL \memory_reg[0][36]  ( .D(n2336), .CP(clk), .Q(\memory[0][36] ) );
  CFD1QXL \memory_reg[0][35]  ( .D(n2337), .CP(clk), .Q(\memory[0][35] ) );
  CFD1QXL \memory_reg[0][34]  ( .D(n2338), .CP(clk), .Q(\memory[0][34] ) );
  CFD1QXL \memory_reg[0][33]  ( .D(n2339), .CP(clk), .Q(\memory[0][33] ) );
  CFD1QXL \memory_reg[0][32]  ( .D(n2340), .CP(clk), .Q(\memory[0][32] ) );
  CFD1QXL \memory_reg[0][31]  ( .D(n2341), .CP(clk), .Q(\memory[0][31] ) );
  CFD1QXL \memory_reg[0][30]  ( .D(n2342), .CP(clk), .Q(\memory[0][30] ) );
  CFD1QXL \memory_reg[0][29]  ( .D(n2343), .CP(clk), .Q(\memory[0][29] ) );
  CFD1QXL \memory_reg[0][28]  ( .D(n2344), .CP(clk), .Q(\memory[0][28] ) );
  CFD1QXL \memory_reg[0][27]  ( .D(n2345), .CP(clk), .Q(\memory[0][27] ) );
  CFD1QXL \memory_reg[0][26]  ( .D(n2346), .CP(clk), .Q(\memory[0][26] ) );
  CFD1QXL \memory_reg[0][25]  ( .D(n2347), .CP(clk), .Q(\memory[0][25] ) );
  CFD1QXL \memory_reg[0][24]  ( .D(n2348), .CP(clk), .Q(\memory[0][24] ) );
  CFD1QXL \memory_reg[0][23]  ( .D(n2349), .CP(clk), .Q(\memory[0][23] ) );
  CFD1QXL \memory_reg[0][22]  ( .D(n2350), .CP(clk), .Q(\memory[0][22] ) );
  CFD1QXL \memory_reg[0][21]  ( .D(n2351), .CP(clk), .Q(\memory[0][21] ) );
  CFD1QXL \memory_reg[0][20]  ( .D(n2352), .CP(clk), .Q(\memory[0][20] ) );
  CFD1QXL \memory_reg[0][19]  ( .D(n2353), .CP(clk), .Q(\memory[0][19] ) );
  CFD1QXL \memory_reg[0][18]  ( .D(n2354), .CP(clk), .Q(\memory[0][18] ) );
  CFD1QXL \memory_reg[0][17]  ( .D(n2355), .CP(clk), .Q(\memory[0][17] ) );
  CFD1QXL \memory_reg[0][16]  ( .D(n2356), .CP(clk), .Q(\memory[0][16] ) );
  CFD1QXL \memory_reg[0][15]  ( .D(n2357), .CP(clk), .Q(\memory[0][15] ) );
  CFD1QXL \memory_reg[0][14]  ( .D(n2358), .CP(clk), .Q(\memory[0][14] ) );
  CFD1QXL \memory_reg[0][13]  ( .D(n2359), .CP(clk), .Q(\memory[0][13] ) );
  CFD1QXL \memory_reg[0][12]  ( .D(n2360), .CP(clk), .Q(\memory[0][12] ) );
  CFD1QXL \memory_reg[0][11]  ( .D(n2361), .CP(clk), .Q(\memory[0][11] ) );
  CFD1QXL \memory_reg[0][10]  ( .D(n2362), .CP(clk), .Q(\memory[0][10] ) );
  CFD1QXL \memory_reg[0][9]  ( .D(n2363), .CP(clk), .Q(\memory[0][9] ) );
  CFD1QXL \memory_reg[0][8]  ( .D(n2364), .CP(clk), .Q(\memory[0][8] ) );
  CFD1QXL \memory_reg[0][7]  ( .D(n2365), .CP(clk), .Q(\memory[0][7] ) );
  CFD1QXL \memory_reg[0][6]  ( .D(n2366), .CP(clk), .Q(\memory[0][6] ) );
  CFD1QXL \memory_reg[0][5]  ( .D(n2367), .CP(clk), .Q(\memory[0][5] ) );
  CFD1QXL \memory_reg[0][4]  ( .D(n2368), .CP(clk), .Q(\memory[0][4] ) );
  CFD1QXL \memory_reg[0][3]  ( .D(n2369), .CP(clk), .Q(\memory[0][3] ) );
  CFD1QXL \memory_reg[0][2]  ( .D(n2370), .CP(clk), .Q(\memory[0][2] ) );
  CFD1QXL \memory_reg[0][1]  ( .D(n2371), .CP(clk), .Q(\memory[0][1] ) );
  CFD1QXL \memory_reg[0][0]  ( .D(n2372), .CP(clk), .Q(\memory[0][0] ) );
  CFD2QX2 \read_ptr_reg[3]  ( .D(n2379), .CP(clk), .CD(n77), .Q(N41) );
  CFD2QX4 \read_ptr_reg[4]  ( .D(n2378), .CP(clk), .CD(n77), .Q(N42) );
  CMX2X2 U2689 ( .A0(counter[3]), .A1(N2536), .S(N4961), .Z(n2456) );
  CMX2X2 U2690 ( .A0(counter[2]), .A1(N2535), .S(N4961), .Z(n2455) );
  CMX2X4 U2691 ( .A0(counter[4]), .A1(N2537), .S(N4961), .Z(n2457) );
  CMX2X2 U2692 ( .A0(counter[1]), .A1(N2534), .S(N4961), .Z(n2454) );
  CMX2X4 U2693 ( .A0(counter[5]), .A1(N2538), .S(N4961), .Z(n2458) );
  CNIVX1 U2694 ( .A(n2460), .Z(n2530) );
  CNIVX1 U2695 ( .A(n2461), .Z(n2531) );
  CNIVX1 U2696 ( .A(n2462), .Z(n2532) );
  CNIVX1 U2697 ( .A(n2463), .Z(n2533) );
  CNIVX1 U2698 ( .A(n2464), .Z(n2534) );
  CNIVX1 U2699 ( .A(n2465), .Z(n2535) );
  CMXI2X2 U2700 ( .A0(n2609), .A1(N115), .S(stopout), .Z(n2608) );
  CMXI2X2 U2701 ( .A0(n2607), .A1(N5117), .S(read), .Z(n2606) );
  CMX2X2 U2702 ( .A0(\memory[31][70] ), .A1(lout_new[6]), .S(N4818), .Z(n101)
         );
  CMX2X2 U2703 ( .A0(\memory[31][69] ), .A1(lout_new[5]), .S(N4818), .Z(n102)
         );
  CMX2X2 U2704 ( .A0(\memory[31][68] ), .A1(lout_new[4]), .S(N4818), .Z(n103)
         );
  CMX2X2 U2705 ( .A0(\memory[31][67] ), .A1(lout_new[3]), .S(N4818), .Z(n104)
         );
  CMX2X2 U2706 ( .A0(\memory[31][66] ), .A1(lout_new[2]), .S(N4818), .Z(n105)
         );
  CMX2X2 U2707 ( .A0(\memory[31][65] ), .A1(lout_new[1]), .S(N4818), .Z(n106)
         );
  CMX2X2 U2708 ( .A0(\memory[31][64] ), .A1(lout_new[0]), .S(N4818), .Z(n107)
         );
  CMX2X2 U2709 ( .A0(\memory[30][70] ), .A1(lout_new[6]), .S(N4747), .Z(n172)
         );
  CMX2X2 U2710 ( .A0(\memory[30][69] ), .A1(lout_new[5]), .S(N4747), .Z(n173)
         );
  CMX2X2 U2711 ( .A0(\memory[30][68] ), .A1(lout_new[4]), .S(N4747), .Z(n174)
         );
  CMX2X2 U2712 ( .A0(\memory[30][67] ), .A1(lout_new[3]), .S(N4747), .Z(n175)
         );
  CMX2X2 U2713 ( .A0(\memory[30][66] ), .A1(lout_new[2]), .S(N4747), .Z(n176)
         );
  CMX2X2 U2714 ( .A0(\memory[30][65] ), .A1(lout_new[1]), .S(N4747), .Z(n177)
         );
  CMX2X2 U2715 ( .A0(\memory[30][64] ), .A1(lout_new[0]), .S(N4747), .Z(n178)
         );
  CMX2X4 U2716 ( .A0(\memory[29][70] ), .A1(lout_new[6]), .S(N4676), .Z(n243)
         );
  CMX2X4 U2717 ( .A0(\memory[29][69] ), .A1(lout_new[5]), .S(N4676), .Z(n244)
         );
  CMX2X4 U2718 ( .A0(\memory[29][68] ), .A1(lout_new[4]), .S(N4676), .Z(n245)
         );
  CMX2X4 U2719 ( .A0(\memory[29][67] ), .A1(lout_new[3]), .S(N4676), .Z(n246)
         );
  CMX2X4 U2720 ( .A0(\memory[29][66] ), .A1(lout_new[2]), .S(N4676), .Z(n247)
         );
  CMX2X4 U2721 ( .A0(\memory[29][65] ), .A1(lout_new[1]), .S(N4676), .Z(n248)
         );
  CMX2X4 U2722 ( .A0(\memory[29][64] ), .A1(lout_new[0]), .S(N4676), .Z(n249)
         );
  CMX2X2 U2723 ( .A0(\memory[28][70] ), .A1(lout_new[6]), .S(N4605), .Z(n314)
         );
  CMX2X2 U2724 ( .A0(\memory[28][69] ), .A1(lout_new[5]), .S(N4605), .Z(n315)
         );
  CMX2X2 U2725 ( .A0(\memory[28][68] ), .A1(lout_new[4]), .S(N4605), .Z(n316)
         );
  CMX2X2 U2726 ( .A0(\memory[28][67] ), .A1(lout_new[3]), .S(N4605), .Z(n317)
         );
  CMX2X2 U2727 ( .A0(\memory[28][66] ), .A1(lout_new[2]), .S(N4605), .Z(n318)
         );
  CMX2X2 U2728 ( .A0(\memory[28][65] ), .A1(lout_new[1]), .S(N4605), .Z(n319)
         );
  CMX2X2 U2729 ( .A0(\memory[28][64] ), .A1(lout_new[0]), .S(N4605), .Z(n320)
         );
  CMX2X2 U2730 ( .A0(\memory[27][70] ), .A1(lout_new[6]), .S(N4534), .Z(n385)
         );
  CMX2X2 U2731 ( .A0(\memory[27][69] ), .A1(lout_new[5]), .S(N4534), .Z(n386)
         );
  CMX2X2 U2732 ( .A0(\memory[27][68] ), .A1(lout_new[4]), .S(N4534), .Z(n387)
         );
  CMX2X2 U2733 ( .A0(\memory[27][67] ), .A1(lout_new[3]), .S(N4534), .Z(n388)
         );
  CMX2X2 U2734 ( .A0(\memory[27][66] ), .A1(lout_new[2]), .S(N4534), .Z(n389)
         );
  CMX2X2 U2735 ( .A0(\memory[27][65] ), .A1(lout_new[1]), .S(N4534), .Z(n390)
         );
  CMX2X2 U2736 ( .A0(\memory[27][64] ), .A1(lout_new[0]), .S(N4534), .Z(n391)
         );
  CMX2X2 U2737 ( .A0(\memory[26][70] ), .A1(lout_new[6]), .S(N4463), .Z(n456)
         );
  CMX2X2 U2738 ( .A0(\memory[26][69] ), .A1(lout_new[5]), .S(N4463), .Z(n457)
         );
  CMX2X2 U2739 ( .A0(\memory[26][68] ), .A1(lout_new[4]), .S(N4463), .Z(n458)
         );
  CMX2X2 U2740 ( .A0(\memory[26][67] ), .A1(lout_new[3]), .S(N4463), .Z(n459)
         );
  CMX2X2 U2741 ( .A0(\memory[26][66] ), .A1(lout_new[2]), .S(N4463), .Z(n460)
         );
  CMX2X2 U2742 ( .A0(\memory[26][65] ), .A1(lout_new[1]), .S(N4463), .Z(n461)
         );
  CMX2X2 U2743 ( .A0(\memory[26][64] ), .A1(lout_new[0]), .S(N4463), .Z(n462)
         );
  CMX2X2 U2744 ( .A0(\memory[25][70] ), .A1(lout_new[6]), .S(N4392), .Z(n527)
         );
  CMX2X2 U2745 ( .A0(\memory[25][69] ), .A1(lout_new[5]), .S(N4392), .Z(n528)
         );
  CMX2X2 U2746 ( .A0(\memory[25][68] ), .A1(lout_new[4]), .S(N4392), .Z(n529)
         );
  CMX2X2 U2747 ( .A0(\memory[25][67] ), .A1(lout_new[3]), .S(N4392), .Z(n530)
         );
  CMX2X2 U2748 ( .A0(\memory[25][66] ), .A1(lout_new[2]), .S(N4392), .Z(n531)
         );
  CMX2X2 U2749 ( .A0(\memory[25][65] ), .A1(lout_new[1]), .S(N4392), .Z(n532)
         );
  CMX2X2 U2750 ( .A0(\memory[25][64] ), .A1(lout_new[0]), .S(N4392), .Z(n533)
         );
  CMX2X2 U2751 ( .A0(\memory[24][70] ), .A1(lout_new[6]), .S(N4321), .Z(n598)
         );
  CMX2X2 U2752 ( .A0(\memory[24][69] ), .A1(lout_new[5]), .S(N4321), .Z(n599)
         );
  CMX2X2 U2753 ( .A0(\memory[24][68] ), .A1(lout_new[4]), .S(N4321), .Z(n600)
         );
  CMX2X2 U2754 ( .A0(\memory[24][67] ), .A1(lout_new[3]), .S(N4321), .Z(n601)
         );
  CMX2X2 U2755 ( .A0(\memory[24][66] ), .A1(lout_new[2]), .S(N4321), .Z(n602)
         );
  CMX2X2 U2756 ( .A0(\memory[24][65] ), .A1(lout_new[1]), .S(N4321), .Z(n603)
         );
  CMX2X2 U2757 ( .A0(\memory[24][64] ), .A1(lout_new[0]), .S(N4321), .Z(n604)
         );
  CMX2X2 U2758 ( .A0(\memory[23][70] ), .A1(lout_new[6]), .S(N4250), .Z(n669)
         );
  CMX2X2 U2759 ( .A0(\memory[23][69] ), .A1(lout_new[5]), .S(N4250), .Z(n670)
         );
  CMX2X2 U2760 ( .A0(\memory[23][68] ), .A1(lout_new[4]), .S(N4250), .Z(n671)
         );
  CMX2X2 U2761 ( .A0(\memory[23][67] ), .A1(lout_new[3]), .S(N4250), .Z(n672)
         );
  CMX2X2 U2762 ( .A0(\memory[23][66] ), .A1(lout_new[2]), .S(N4250), .Z(n673)
         );
  CMX2X2 U2763 ( .A0(\memory[23][65] ), .A1(lout_new[1]), .S(N4250), .Z(n674)
         );
  CMX2X2 U2764 ( .A0(\memory[23][64] ), .A1(lout_new[0]), .S(N4250), .Z(n675)
         );
  CMX2X2 U2765 ( .A0(\memory[22][70] ), .A1(lout_new[6]), .S(N4179), .Z(n740)
         );
  CMX2X2 U2766 ( .A0(\memory[22][69] ), .A1(lout_new[5]), .S(N4179), .Z(n741)
         );
  CMX2X2 U2767 ( .A0(\memory[22][68] ), .A1(lout_new[4]), .S(N4179), .Z(n742)
         );
  CMX2X2 U2768 ( .A0(\memory[22][67] ), .A1(lout_new[3]), .S(N4179), .Z(n743)
         );
  CMX2X2 U2769 ( .A0(\memory[22][66] ), .A1(lout_new[2]), .S(N4179), .Z(n744)
         );
  CMX2X2 U2770 ( .A0(\memory[22][65] ), .A1(lout_new[1]), .S(N4179), .Z(n745)
         );
  CMX2X2 U2771 ( .A0(\memory[22][64] ), .A1(lout_new[0]), .S(N4179), .Z(n746)
         );
  CMX2X4 U2772 ( .A0(\memory[21][70] ), .A1(lout_new[6]), .S(N4108), .Z(n811)
         );
  CMX2X4 U2773 ( .A0(\memory[21][69] ), .A1(lout_new[5]), .S(N4108), .Z(n812)
         );
  CMX2X4 U2774 ( .A0(\memory[21][68] ), .A1(lout_new[4]), .S(N4108), .Z(n813)
         );
  CMX2X4 U2775 ( .A0(\memory[21][67] ), .A1(lout_new[3]), .S(N4108), .Z(n814)
         );
  CMX2X4 U2776 ( .A0(\memory[21][66] ), .A1(lout_new[2]), .S(N4108), .Z(n815)
         );
  CMX2X4 U2777 ( .A0(\memory[21][65] ), .A1(lout_new[1]), .S(N4108), .Z(n816)
         );
  CMX2X4 U2778 ( .A0(\memory[21][64] ), .A1(lout_new[0]), .S(N4108), .Z(n817)
         );
  CMX2X2 U2779 ( .A0(\memory[20][70] ), .A1(lout_new[6]), .S(N4037), .Z(n882)
         );
  CMX2X2 U2780 ( .A0(\memory[20][69] ), .A1(lout_new[5]), .S(N4037), .Z(n883)
         );
  CMX2X2 U2781 ( .A0(\memory[20][68] ), .A1(lout_new[4]), .S(N4037), .Z(n884)
         );
  CMX2X2 U2782 ( .A0(\memory[20][67] ), .A1(lout_new[3]), .S(N4037), .Z(n885)
         );
  CMX2X2 U2783 ( .A0(\memory[20][66] ), .A1(lout_new[2]), .S(N4037), .Z(n886)
         );
  CMX2X2 U2784 ( .A0(\memory[20][65] ), .A1(lout_new[1]), .S(N4037), .Z(n887)
         );
  CMX2X2 U2785 ( .A0(\memory[20][64] ), .A1(lout_new[0]), .S(N4037), .Z(n888)
         );
  CMX2X2 U2786 ( .A0(\memory[19][70] ), .A1(lout_new[6]), .S(N3966), .Z(n953)
         );
  CMX2X2 U2787 ( .A0(\memory[19][69] ), .A1(lout_new[5]), .S(N3966), .Z(n954)
         );
  CMX2X2 U2788 ( .A0(\memory[19][68] ), .A1(lout_new[4]), .S(N3966), .Z(n955)
         );
  CMX2X2 U2789 ( .A0(\memory[19][67] ), .A1(lout_new[3]), .S(N3966), .Z(n956)
         );
  CMX2X2 U2790 ( .A0(\memory[19][66] ), .A1(lout_new[2]), .S(N3966), .Z(n957)
         );
  CMX2X2 U2791 ( .A0(\memory[19][65] ), .A1(lout_new[1]), .S(N3966), .Z(n958)
         );
  CMX2X2 U2792 ( .A0(\memory[19][64] ), .A1(lout_new[0]), .S(N3966), .Z(n959)
         );
  CMX2X2 U2793 ( .A0(\memory[18][70] ), .A1(lout_new[6]), .S(N3895), .Z(n1024)
         );
  CMX2X2 U2794 ( .A0(\memory[18][69] ), .A1(lout_new[5]), .S(N3895), .Z(n1025)
         );
  CMX2X2 U2795 ( .A0(\memory[18][68] ), .A1(lout_new[4]), .S(N3895), .Z(n1026)
         );
  CMX2X2 U2796 ( .A0(\memory[18][67] ), .A1(lout_new[3]), .S(N3895), .Z(n1027)
         );
  CMX2X2 U2797 ( .A0(\memory[18][66] ), .A1(lout_new[2]), .S(N3895), .Z(n1028)
         );
  CMX2X2 U2798 ( .A0(\memory[18][65] ), .A1(lout_new[1]), .S(N3895), .Z(n1029)
         );
  CMX2X2 U2799 ( .A0(\memory[18][64] ), .A1(lout_new[0]), .S(N3895), .Z(n1030)
         );
  CMX2X2 U2800 ( .A0(\memory[17][70] ), .A1(lout_new[6]), .S(N3824), .Z(n1095)
         );
  CMX2X2 U2801 ( .A0(\memory[17][69] ), .A1(lout_new[5]), .S(N3824), .Z(n1096)
         );
  CMX2X2 U2802 ( .A0(\memory[17][68] ), .A1(lout_new[4]), .S(N3824), .Z(n1097)
         );
  CMX2X2 U2803 ( .A0(\memory[17][67] ), .A1(lout_new[3]), .S(N3824), .Z(n1098)
         );
  CMX2X2 U2804 ( .A0(\memory[17][66] ), .A1(lout_new[2]), .S(N3824), .Z(n1099)
         );
  CMX2X2 U2805 ( .A0(\memory[17][65] ), .A1(lout_new[1]), .S(N3824), .Z(n1100)
         );
  CMX2X2 U2806 ( .A0(\memory[17][64] ), .A1(lout_new[0]), .S(N3824), .Z(n1101)
         );
  CMX2X2 U2807 ( .A0(\memory[16][70] ), .A1(lout_new[6]), .S(N3753), .Z(n1166)
         );
  CMX2X2 U2808 ( .A0(\memory[16][69] ), .A1(lout_new[5]), .S(N3753), .Z(n1167)
         );
  CMX2X2 U2809 ( .A0(\memory[16][68] ), .A1(lout_new[4]), .S(N3753), .Z(n1168)
         );
  CMX2X2 U2810 ( .A0(\memory[16][67] ), .A1(lout_new[3]), .S(N3753), .Z(n1169)
         );
  CMX2X2 U2811 ( .A0(\memory[16][66] ), .A1(lout_new[2]), .S(N3753), .Z(n1170)
         );
  CMX2X2 U2812 ( .A0(\memory[16][65] ), .A1(lout_new[1]), .S(N3753), .Z(n1171)
         );
  CMX2X2 U2813 ( .A0(\memory[16][64] ), .A1(lout_new[0]), .S(N3753), .Z(n1172)
         );
  CMX2X2 U2814 ( .A0(\memory[15][70] ), .A1(lout_new[6]), .S(N3682), .Z(n1237)
         );
  CMX2X2 U2815 ( .A0(\memory[15][69] ), .A1(lout_new[5]), .S(N3682), .Z(n1238)
         );
  CMX2X2 U2816 ( .A0(\memory[15][68] ), .A1(lout_new[4]), .S(N3682), .Z(n1239)
         );
  CMX2X2 U2817 ( .A0(\memory[15][67] ), .A1(lout_new[3]), .S(N3682), .Z(n1240)
         );
  CMX2X2 U2818 ( .A0(\memory[15][66] ), .A1(lout_new[2]), .S(N3682), .Z(n1241)
         );
  CMX2X2 U2819 ( .A0(\memory[15][65] ), .A1(lout_new[1]), .S(N3682), .Z(n1242)
         );
  CMX2X2 U2820 ( .A0(\memory[15][64] ), .A1(lout_new[0]), .S(N3682), .Z(n1243)
         );
  CMX2X2 U2821 ( .A0(\memory[14][70] ), .A1(lout_new[6]), .S(N3611), .Z(n1308)
         );
  CMX2X2 U2822 ( .A0(\memory[14][69] ), .A1(lout_new[5]), .S(N3611), .Z(n1309)
         );
  CMX2X2 U2823 ( .A0(\memory[14][68] ), .A1(lout_new[4]), .S(N3611), .Z(n1310)
         );
  CMX2X2 U2824 ( .A0(\memory[14][67] ), .A1(lout_new[3]), .S(N3611), .Z(n1311)
         );
  CMX2X2 U2825 ( .A0(\memory[14][66] ), .A1(lout_new[2]), .S(N3611), .Z(n1312)
         );
  CMX2X2 U2826 ( .A0(\memory[14][65] ), .A1(lout_new[1]), .S(N3611), .Z(n1313)
         );
  CMX2X2 U2827 ( .A0(\memory[14][64] ), .A1(lout_new[0]), .S(N3611), .Z(n1314)
         );
  CMX2X4 U2828 ( .A0(\memory[13][70] ), .A1(lout_new[6]), .S(N3540), .Z(n1379)
         );
  CMX2X4 U2829 ( .A0(\memory[13][69] ), .A1(lout_new[5]), .S(N3540), .Z(n1380)
         );
  CMX2X4 U2830 ( .A0(\memory[13][68] ), .A1(lout_new[4]), .S(N3540), .Z(n1381)
         );
  CMX2X4 U2831 ( .A0(\memory[13][67] ), .A1(lout_new[3]), .S(N3540), .Z(n1382)
         );
  CMX2X4 U2832 ( .A0(\memory[13][66] ), .A1(lout_new[2]), .S(N3540), .Z(n1383)
         );
  CMX2X4 U2833 ( .A0(\memory[13][65] ), .A1(lout_new[1]), .S(N3540), .Z(n1384)
         );
  CMX2X4 U2834 ( .A0(\memory[13][64] ), .A1(lout_new[0]), .S(N3540), .Z(n1385)
         );
  CMX2X2 U2835 ( .A0(\memory[12][70] ), .A1(lout_new[6]), .S(N3469), .Z(n1450)
         );
  CMX2X2 U2836 ( .A0(\memory[12][69] ), .A1(lout_new[5]), .S(N3469), .Z(n1451)
         );
  CMX2X2 U2837 ( .A0(\memory[12][68] ), .A1(lout_new[4]), .S(N3469), .Z(n1452)
         );
  CMX2X2 U2838 ( .A0(\memory[12][67] ), .A1(lout_new[3]), .S(N3469), .Z(n1453)
         );
  CMX2X2 U2839 ( .A0(\memory[12][66] ), .A1(lout_new[2]), .S(N3469), .Z(n1454)
         );
  CMX2X2 U2840 ( .A0(\memory[12][65] ), .A1(lout_new[1]), .S(N3469), .Z(n1455)
         );
  CMX2X2 U2841 ( .A0(\memory[12][64] ), .A1(lout_new[0]), .S(N3469), .Z(n1456)
         );
  CMX2X2 U2842 ( .A0(\memory[11][70] ), .A1(lout_new[6]), .S(N3398), .Z(n1521)
         );
  CMX2X2 U2843 ( .A0(\memory[11][69] ), .A1(lout_new[5]), .S(N3398), .Z(n1522)
         );
  CMX2X2 U2844 ( .A0(\memory[11][68] ), .A1(lout_new[4]), .S(N3398), .Z(n1523)
         );
  CMX2X2 U2845 ( .A0(\memory[11][67] ), .A1(lout_new[3]), .S(N3398), .Z(n1524)
         );
  CMX2X2 U2846 ( .A0(\memory[11][66] ), .A1(lout_new[2]), .S(N3398), .Z(n1525)
         );
  CMX2X2 U2847 ( .A0(\memory[11][65] ), .A1(lout_new[1]), .S(N3398), .Z(n1526)
         );
  CMX2X2 U2848 ( .A0(\memory[11][64] ), .A1(lout_new[0]), .S(N3398), .Z(n1527)
         );
  CMX2X2 U2849 ( .A0(\memory[10][70] ), .A1(lout_new[6]), .S(N3327), .Z(n1592)
         );
  CMX2X2 U2850 ( .A0(\memory[10][69] ), .A1(lout_new[5]), .S(N3327), .Z(n1593)
         );
  CMX2X2 U2851 ( .A0(\memory[10][68] ), .A1(lout_new[4]), .S(N3327), .Z(n1594)
         );
  CMX2X2 U2852 ( .A0(\memory[10][67] ), .A1(lout_new[3]), .S(N3327), .Z(n1595)
         );
  CMX2X2 U2853 ( .A0(\memory[10][66] ), .A1(lout_new[2]), .S(N3327), .Z(n1596)
         );
  CMX2X2 U2854 ( .A0(\memory[10][65] ), .A1(lout_new[1]), .S(N3327), .Z(n1597)
         );
  CMX2X2 U2855 ( .A0(\memory[10][64] ), .A1(lout_new[0]), .S(N3327), .Z(n1598)
         );
  CMX2X2 U2856 ( .A0(\memory[9][70] ), .A1(lout_new[6]), .S(N3256), .Z(n1663)
         );
  CMX2X2 U2857 ( .A0(\memory[9][69] ), .A1(lout_new[5]), .S(N3256), .Z(n1664)
         );
  CMX2X2 U2858 ( .A0(\memory[9][68] ), .A1(lout_new[4]), .S(N3256), .Z(n1665)
         );
  CMX2X2 U2859 ( .A0(\memory[9][67] ), .A1(lout_new[3]), .S(N3256), .Z(n1666)
         );
  CMX2X2 U2860 ( .A0(\memory[9][66] ), .A1(lout_new[2]), .S(N3256), .Z(n1667)
         );
  CMX2X2 U2861 ( .A0(\memory[9][65] ), .A1(lout_new[1]), .S(N3256), .Z(n1668)
         );
  CMX2X2 U2862 ( .A0(\memory[9][64] ), .A1(lout_new[0]), .S(N3256), .Z(n1669)
         );
  CMX2X2 U2863 ( .A0(\memory[8][70] ), .A1(lout_new[6]), .S(N3185), .Z(n1734)
         );
  CMX2X2 U2864 ( .A0(\memory[8][69] ), .A1(lout_new[5]), .S(N3185), .Z(n1735)
         );
  CMX2X2 U2865 ( .A0(\memory[8][68] ), .A1(lout_new[4]), .S(N3185), .Z(n1736)
         );
  CMX2X2 U2866 ( .A0(\memory[8][67] ), .A1(lout_new[3]), .S(N3185), .Z(n1737)
         );
  CMX2X2 U2867 ( .A0(\memory[8][66] ), .A1(lout_new[2]), .S(N3185), .Z(n1738)
         );
  CMX2X2 U2868 ( .A0(\memory[8][65] ), .A1(lout_new[1]), .S(N3185), .Z(n1739)
         );
  CMX2X2 U2869 ( .A0(\memory[8][64] ), .A1(lout_new[0]), .S(N3185), .Z(n1740)
         );
  CMX2X2 U2870 ( .A0(\memory[7][70] ), .A1(lout_new[6]), .S(N3114), .Z(n1805)
         );
  CMX2X2 U2871 ( .A0(\memory[7][69] ), .A1(lout_new[5]), .S(N3114), .Z(n1806)
         );
  CMX2X2 U2872 ( .A0(\memory[7][68] ), .A1(lout_new[4]), .S(N3114), .Z(n1807)
         );
  CMX2X2 U2873 ( .A0(\memory[7][67] ), .A1(lout_new[3]), .S(N3114), .Z(n1808)
         );
  CMX2X2 U2874 ( .A0(\memory[7][66] ), .A1(lout_new[2]), .S(N3114), .Z(n1809)
         );
  CMX2X2 U2875 ( .A0(\memory[7][65] ), .A1(lout_new[1]), .S(N3114), .Z(n1810)
         );
  CMX2X2 U2876 ( .A0(\memory[7][64] ), .A1(lout_new[0]), .S(N3114), .Z(n1811)
         );
  CMX2X2 U2877 ( .A0(\memory[6][70] ), .A1(lout_new[6]), .S(N3043), .Z(n1876)
         );
  CMX2X2 U2878 ( .A0(\memory[6][69] ), .A1(lout_new[5]), .S(N3043), .Z(n1877)
         );
  CMX2X2 U2879 ( .A0(\memory[6][68] ), .A1(lout_new[4]), .S(N3043), .Z(n1878)
         );
  CMX2X2 U2880 ( .A0(\memory[6][67] ), .A1(lout_new[3]), .S(N3043), .Z(n1879)
         );
  CMX2X2 U2881 ( .A0(\memory[6][66] ), .A1(lout_new[2]), .S(N3043), .Z(n1880)
         );
  CMX2X2 U2882 ( .A0(\memory[6][65] ), .A1(lout_new[1]), .S(N3043), .Z(n1881)
         );
  CMX2X2 U2883 ( .A0(\memory[6][64] ), .A1(lout_new[0]), .S(N3043), .Z(n1882)
         );
  CMX2X4 U2884 ( .A0(\memory[5][70] ), .A1(lout_new[6]), .S(N2972), .Z(n1947)
         );
  CMX2X4 U2885 ( .A0(\memory[5][69] ), .A1(lout_new[5]), .S(N2972), .Z(n1948)
         );
  CMX2X4 U2886 ( .A0(\memory[5][68] ), .A1(lout_new[4]), .S(N2972), .Z(n1949)
         );
  CMX2X4 U2887 ( .A0(\memory[5][67] ), .A1(lout_new[3]), .S(N2972), .Z(n1950)
         );
  CMX2X4 U2888 ( .A0(\memory[5][66] ), .A1(lout_new[2]), .S(N2972), .Z(n1951)
         );
  CMX2X4 U2889 ( .A0(\memory[5][65] ), .A1(lout_new[1]), .S(N2972), .Z(n1952)
         );
  CMX2X4 U2890 ( .A0(\memory[5][64] ), .A1(lout_new[0]), .S(N2972), .Z(n1953)
         );
  CMX2X2 U2891 ( .A0(\memory[4][70] ), .A1(lout_new[6]), .S(N2901), .Z(n2018)
         );
  CMX2X2 U2892 ( .A0(\memory[4][69] ), .A1(lout_new[5]), .S(N2901), .Z(n2019)
         );
  CMX2X2 U2893 ( .A0(\memory[4][68] ), .A1(lout_new[4]), .S(N2901), .Z(n2020)
         );
  CMX2X2 U2894 ( .A0(\memory[4][67] ), .A1(lout_new[3]), .S(N2901), .Z(n2021)
         );
  CMX2X2 U2895 ( .A0(\memory[4][66] ), .A1(lout_new[2]), .S(N2901), .Z(n2022)
         );
  CMX2X2 U2896 ( .A0(\memory[4][65] ), .A1(lout_new[1]), .S(N2901), .Z(n2023)
         );
  CMX2X2 U2897 ( .A0(\memory[4][64] ), .A1(lout_new[0]), .S(N2901), .Z(n2024)
         );
  CMX2X2 U2898 ( .A0(\memory[3][70] ), .A1(lout_new[6]), .S(N2830), .Z(n2089)
         );
  CMX2X2 U2899 ( .A0(\memory[3][69] ), .A1(lout_new[5]), .S(N2830), .Z(n2090)
         );
  CMX2X2 U2900 ( .A0(\memory[3][68] ), .A1(lout_new[4]), .S(N2830), .Z(n2091)
         );
  CMX2X2 U2901 ( .A0(\memory[3][67] ), .A1(lout_new[3]), .S(N2830), .Z(n2092)
         );
  CMX2X2 U2902 ( .A0(\memory[3][66] ), .A1(lout_new[2]), .S(N2830), .Z(n2093)
         );
  CMX2X2 U2903 ( .A0(\memory[3][65] ), .A1(lout_new[1]), .S(N2830), .Z(n2094)
         );
  CMX2X2 U2904 ( .A0(\memory[3][64] ), .A1(lout_new[0]), .S(N2830), .Z(n2095)
         );
  CMX2X2 U2905 ( .A0(\memory[2][70] ), .A1(lout_new[6]), .S(N2759), .Z(n2160)
         );
  CMX2X2 U2906 ( .A0(\memory[2][69] ), .A1(lout_new[5]), .S(N2759), .Z(n2161)
         );
  CMX2X2 U2907 ( .A0(\memory[2][68] ), .A1(lout_new[4]), .S(N2759), .Z(n2162)
         );
  CMX2X2 U2908 ( .A0(\memory[2][67] ), .A1(lout_new[3]), .S(N2759), .Z(n2163)
         );
  CMX2X2 U2909 ( .A0(\memory[2][66] ), .A1(lout_new[2]), .S(N2759), .Z(n2164)
         );
  CMX2X2 U2910 ( .A0(\memory[2][65] ), .A1(lout_new[1]), .S(N2759), .Z(n2165)
         );
  CMX2X2 U2911 ( .A0(\memory[2][64] ), .A1(lout_new[0]), .S(N2759), .Z(n2166)
         );
  CMX2X2 U2912 ( .A0(\memory[1][70] ), .A1(lout_new[6]), .S(N2688), .Z(n2231)
         );
  CMX2X2 U2913 ( .A0(\memory[1][69] ), .A1(lout_new[5]), .S(N2688), .Z(n2232)
         );
  CMX2X2 U2914 ( .A0(\memory[1][68] ), .A1(lout_new[4]), .S(N2688), .Z(n2233)
         );
  CMX2X2 U2915 ( .A0(\memory[1][67] ), .A1(lout_new[3]), .S(N2688), .Z(n2234)
         );
  CMX2X2 U2916 ( .A0(\memory[1][66] ), .A1(lout_new[2]), .S(N2688), .Z(n2235)
         );
  CMX2X2 U2917 ( .A0(\memory[1][65] ), .A1(lout_new[1]), .S(N2688), .Z(n2236)
         );
  CMX2X2 U2918 ( .A0(\memory[1][64] ), .A1(lout_new[0]), .S(N2688), .Z(n2237)
         );
  CMX2X2 U2919 ( .A0(\memory[0][70] ), .A1(lout_new[6]), .S(N2617), .Z(n2302)
         );
  CMX2X2 U2920 ( .A0(\memory[0][69] ), .A1(lout_new[5]), .S(N2617), .Z(n2303)
         );
  CMX2X2 U2921 ( .A0(\memory[0][68] ), .A1(lout_new[4]), .S(N2617), .Z(n2304)
         );
  CMX2X2 U2922 ( .A0(\memory[0][67] ), .A1(lout_new[3]), .S(N2617), .Z(n2305)
         );
  CMX2X2 U2923 ( .A0(\memory[0][66] ), .A1(lout_new[2]), .S(N2617), .Z(n2306)
         );
  CMX2X2 U2924 ( .A0(\memory[0][65] ), .A1(lout_new[1]), .S(N2617), .Z(n2307)
         );
  CMX2X2 U2925 ( .A0(\memory[0][64] ), .A1(lout_new[0]), .S(N2617), .Z(n2308)
         );
  CMX2X2 U2926 ( .A0(\memory[31][63] ), .A1(out_new[63]), .S(N4811), .Z(n108)
         );
  CMX2X2 U2927 ( .A0(\memory[31][62] ), .A1(out_new[62]), .S(N4811), .Z(n109)
         );
  CMX2X2 U2928 ( .A0(\memory[31][61] ), .A1(out_new[61]), .S(N4811), .Z(n110)
         );
  CMX2X2 U2929 ( .A0(\memory[31][60] ), .A1(out_new[60]), .S(N4811), .Z(n111)
         );
  CMX2X2 U2930 ( .A0(\memory[31][59] ), .A1(out_new[59]), .S(N4811), .Z(n112)
         );
  CMX2X2 U2931 ( .A0(\memory[31][58] ), .A1(out_new[58]), .S(N4811), .Z(n113)
         );
  CMX2X2 U2932 ( .A0(\memory[31][57] ), .A1(out_new[57]), .S(N4811), .Z(n114)
         );
  CMX2X2 U2933 ( .A0(\memory[31][56] ), .A1(out_new[56]), .S(N4811), .Z(n115)
         );
  CMX2X2 U2934 ( .A0(\memory[31][55] ), .A1(out_new[55]), .S(N4811), .Z(n116)
         );
  CMX2X2 U2935 ( .A0(\memory[31][54] ), .A1(out_new[54]), .S(N4811), .Z(n117)
         );
  CMX2X2 U2936 ( .A0(\memory[31][53] ), .A1(out_new[53]), .S(N4811), .Z(n118)
         );
  CMX2X2 U2937 ( .A0(\memory[31][52] ), .A1(out_new[52]), .S(N4811), .Z(n119)
         );
  CMX2X2 U2938 ( .A0(\memory[31][51] ), .A1(out_new[51]), .S(N4811), .Z(n120)
         );
  CMX2X2 U2939 ( .A0(\memory[31][50] ), .A1(out_new[50]), .S(N4811), .Z(n121)
         );
  CMX2X2 U2940 ( .A0(\memory[31][49] ), .A1(out_new[49]), .S(N4811), .Z(n122)
         );
  CMX2X2 U2941 ( .A0(\memory[31][48] ), .A1(out_new[48]), .S(N4811), .Z(n123)
         );
  CMX2X2 U2942 ( .A0(\memory[31][47] ), .A1(out_new[47]), .S(N4811), .Z(n124)
         );
  CMX2X2 U2943 ( .A0(\memory[31][46] ), .A1(out_new[46]), .S(N4811), .Z(n125)
         );
  CMX2X2 U2944 ( .A0(\memory[31][45] ), .A1(out_new[45]), .S(N4811), .Z(n126)
         );
  CMX2X2 U2945 ( .A0(\memory[31][44] ), .A1(out_new[44]), .S(N4811), .Z(n127)
         );
  CMX2X2 U2946 ( .A0(\memory[31][43] ), .A1(out_new[43]), .S(N4811), .Z(n128)
         );
  CMX2X2 U2947 ( .A0(\memory[31][42] ), .A1(out_new[42]), .S(N4811), .Z(n129)
         );
  CMX2X2 U2948 ( .A0(\memory[31][41] ), .A1(out_new[41]), .S(N4811), .Z(n130)
         );
  CMX2X2 U2949 ( .A0(\memory[31][40] ), .A1(out_new[40]), .S(N4811), .Z(n131)
         );
  CMX2X2 U2950 ( .A0(\memory[31][39] ), .A1(out_new[39]), .S(N4811), .Z(n132)
         );
  CMX2X2 U2951 ( .A0(\memory[31][38] ), .A1(out_new[38]), .S(N4811), .Z(n133)
         );
  CMX2X2 U2952 ( .A0(\memory[31][37] ), .A1(out_new[37]), .S(N4811), .Z(n134)
         );
  CMX2X2 U2953 ( .A0(\memory[31][36] ), .A1(out_new[36]), .S(N4811), .Z(n135)
         );
  CMX2X2 U2954 ( .A0(\memory[31][35] ), .A1(out_new[35]), .S(N4811), .Z(n136)
         );
  CMX2X2 U2955 ( .A0(\memory[31][34] ), .A1(out_new[34]), .S(N4811), .Z(n137)
         );
  CMX2X2 U2956 ( .A0(\memory[31][33] ), .A1(out_new[33]), .S(N4811), .Z(n138)
         );
  CMX2X2 U2957 ( .A0(\memory[31][32] ), .A1(out_new[32]), .S(N4811), .Z(n139)
         );
  CMX2X2 U2958 ( .A0(\memory[31][31] ), .A1(out_new[31]), .S(N4811), .Z(n140)
         );
  CMX2X2 U2959 ( .A0(\memory[31][30] ), .A1(out_new[30]), .S(N4811), .Z(n141)
         );
  CMX2X2 U2960 ( .A0(\memory[31][29] ), .A1(out_new[29]), .S(N4811), .Z(n142)
         );
  CMX2X2 U2961 ( .A0(\memory[31][28] ), .A1(out_new[28]), .S(N4811), .Z(n143)
         );
  CMX2X2 U2962 ( .A0(\memory[31][27] ), .A1(out_new[27]), .S(N4811), .Z(n144)
         );
  CMX2X2 U2963 ( .A0(\memory[31][26] ), .A1(out_new[26]), .S(N4811), .Z(n145)
         );
  CMX2X2 U2964 ( .A0(\memory[31][25] ), .A1(out_new[25]), .S(N4811), .Z(n146)
         );
  CMX2X2 U2965 ( .A0(\memory[31][24] ), .A1(out_new[24]), .S(N4811), .Z(n147)
         );
  CMX2X2 U2966 ( .A0(\memory[31][23] ), .A1(out_new[23]), .S(N4811), .Z(n148)
         );
  CMX2X2 U2967 ( .A0(\memory[31][22] ), .A1(out_new[22]), .S(N4811), .Z(n149)
         );
  CMX2X2 U2968 ( .A0(\memory[31][21] ), .A1(out_new[21]), .S(N4811), .Z(n150)
         );
  CMX2X2 U2969 ( .A0(\memory[31][20] ), .A1(out_new[20]), .S(N4811), .Z(n151)
         );
  CMX2X2 U2970 ( .A0(\memory[31][19] ), .A1(out_new[19]), .S(N4811), .Z(n152)
         );
  CMX2X2 U2971 ( .A0(\memory[31][18] ), .A1(out_new[18]), .S(N4811), .Z(n153)
         );
  CMX2X2 U2972 ( .A0(\memory[31][17] ), .A1(out_new[17]), .S(N4811), .Z(n154)
         );
  CMX2X2 U2973 ( .A0(\memory[31][16] ), .A1(out_new[16]), .S(N4811), .Z(n155)
         );
  CMX2X2 U2974 ( .A0(\memory[31][15] ), .A1(out_new[15]), .S(N4811), .Z(n156)
         );
  CMX2X2 U2975 ( .A0(\memory[31][14] ), .A1(out_new[14]), .S(N4811), .Z(n157)
         );
  CMX2X2 U2976 ( .A0(\memory[31][13] ), .A1(out_new[13]), .S(N4811), .Z(n158)
         );
  CMX2X2 U2977 ( .A0(\memory[31][12] ), .A1(out_new[12]), .S(N4811), .Z(n159)
         );
  CMX2X2 U2978 ( .A0(\memory[31][11] ), .A1(out_new[11]), .S(N4811), .Z(n160)
         );
  CMX2X2 U2979 ( .A0(\memory[31][10] ), .A1(out_new[10]), .S(N4811), .Z(n161)
         );
  CMX2X2 U2980 ( .A0(\memory[31][9] ), .A1(out_new[9]), .S(N4811), .Z(n162) );
  CMX2X2 U2981 ( .A0(\memory[31][8] ), .A1(out_new[8]), .S(N4811), .Z(n163) );
  CMX2X2 U2982 ( .A0(\memory[31][7] ), .A1(out_new[7]), .S(N4811), .Z(n164) );
  CMX2X2 U2983 ( .A0(\memory[31][6] ), .A1(out_new[6]), .S(N4811), .Z(n165) );
  CMX2X2 U2984 ( .A0(\memory[31][5] ), .A1(out_new[5]), .S(N4811), .Z(n166) );
  CMX2X2 U2985 ( .A0(\memory[31][4] ), .A1(out_new[4]), .S(N4811), .Z(n167) );
  CMX2X2 U2986 ( .A0(\memory[31][3] ), .A1(out_new[3]), .S(N4811), .Z(n168) );
  CMX2X2 U2987 ( .A0(\memory[31][2] ), .A1(out_new[2]), .S(N4811), .Z(n169) );
  CMX2X2 U2988 ( .A0(\memory[31][1] ), .A1(out_new[1]), .S(N4811), .Z(n170) );
  CMX2X2 U2989 ( .A0(\memory[31][0] ), .A1(out_new[0]), .S(N4811), .Z(n171) );
  CMX2X2 U2990 ( .A0(\memory[7][63] ), .A1(out_new[63]), .S(N3107), .Z(n1812)
         );
  CMX2X2 U2991 ( .A0(\memory[7][62] ), .A1(out_new[62]), .S(N3107), .Z(n1813)
         );
  CMX2X2 U2992 ( .A0(\memory[7][61] ), .A1(out_new[61]), .S(N3107), .Z(n1814)
         );
  CMX2X2 U2993 ( .A0(\memory[7][60] ), .A1(out_new[60]), .S(N3107), .Z(n1815)
         );
  CMX2X2 U2994 ( .A0(\memory[7][59] ), .A1(out_new[59]), .S(N3107), .Z(n1816)
         );
  CMX2X2 U2995 ( .A0(\memory[7][58] ), .A1(out_new[58]), .S(N3107), .Z(n1817)
         );
  CMX2X2 U2996 ( .A0(\memory[7][57] ), .A1(out_new[57]), .S(N3107), .Z(n1818)
         );
  CMX2X2 U2997 ( .A0(\memory[7][56] ), .A1(out_new[56]), .S(N3107), .Z(n1819)
         );
  CMX2X2 U2998 ( .A0(\memory[7][55] ), .A1(out_new[55]), .S(N3107), .Z(n1820)
         );
  CMX2X2 U2999 ( .A0(\memory[7][54] ), .A1(out_new[54]), .S(N3107), .Z(n1821)
         );
  CMX2X2 U3000 ( .A0(\memory[7][53] ), .A1(out_new[53]), .S(N3107), .Z(n1822)
         );
  CMX2X2 U3001 ( .A0(\memory[7][52] ), .A1(out_new[52]), .S(N3107), .Z(n1823)
         );
  CMX2X2 U3002 ( .A0(\memory[7][51] ), .A1(out_new[51]), .S(N3107), .Z(n1824)
         );
  CMX2X2 U3003 ( .A0(\memory[7][50] ), .A1(out_new[50]), .S(N3107), .Z(n1825)
         );
  CMX2X2 U3004 ( .A0(\memory[7][49] ), .A1(out_new[49]), .S(N3107), .Z(n1826)
         );
  CMX2X2 U3005 ( .A0(\memory[7][48] ), .A1(out_new[48]), .S(N3107), .Z(n1827)
         );
  CMX2X2 U3006 ( .A0(\memory[7][47] ), .A1(out_new[47]), .S(N3107), .Z(n1828)
         );
  CMX2X2 U3007 ( .A0(\memory[7][46] ), .A1(out_new[46]), .S(N3107), .Z(n1829)
         );
  CMX2X2 U3008 ( .A0(\memory[7][45] ), .A1(out_new[45]), .S(N3107), .Z(n1830)
         );
  CMX2X2 U3009 ( .A0(\memory[7][44] ), .A1(out_new[44]), .S(N3107), .Z(n1831)
         );
  CMX2X2 U3010 ( .A0(\memory[7][43] ), .A1(out_new[43]), .S(N3107), .Z(n1832)
         );
  CMX2X2 U3011 ( .A0(\memory[7][42] ), .A1(out_new[42]), .S(N3107), .Z(n1833)
         );
  CMX2X2 U3012 ( .A0(\memory[7][41] ), .A1(out_new[41]), .S(N3107), .Z(n1834)
         );
  CMX2X2 U3013 ( .A0(\memory[7][40] ), .A1(out_new[40]), .S(N3107), .Z(n1835)
         );
  CMX2X2 U3014 ( .A0(\memory[7][39] ), .A1(out_new[39]), .S(N3107), .Z(n1836)
         );
  CMX2X2 U3015 ( .A0(\memory[7][38] ), .A1(out_new[38]), .S(N3107), .Z(n1837)
         );
  CMX2X2 U3016 ( .A0(\memory[7][37] ), .A1(out_new[37]), .S(N3107), .Z(n1838)
         );
  CMX2X2 U3017 ( .A0(\memory[7][36] ), .A1(out_new[36]), .S(N3107), .Z(n1839)
         );
  CMX2X2 U3018 ( .A0(\memory[7][35] ), .A1(out_new[35]), .S(N3107), .Z(n1840)
         );
  CMX2X2 U3019 ( .A0(\memory[7][34] ), .A1(out_new[34]), .S(N3107), .Z(n1841)
         );
  CMX2X2 U3020 ( .A0(\memory[7][33] ), .A1(out_new[33]), .S(N3107), .Z(n1842)
         );
  CMX2X2 U3021 ( .A0(\memory[7][32] ), .A1(out_new[32]), .S(N3107), .Z(n1843)
         );
  CMX2X2 U3022 ( .A0(\memory[7][31] ), .A1(out_new[31]), .S(N3107), .Z(n1844)
         );
  CMX2X2 U3023 ( .A0(\memory[7][30] ), .A1(out_new[30]), .S(N3107), .Z(n1845)
         );
  CMX2X2 U3024 ( .A0(\memory[7][29] ), .A1(out_new[29]), .S(N3107), .Z(n1846)
         );
  CMX2X2 U3025 ( .A0(\memory[7][28] ), .A1(out_new[28]), .S(N3107), .Z(n1847)
         );
  CMX2X2 U3026 ( .A0(\memory[7][27] ), .A1(out_new[27]), .S(N3107), .Z(n1848)
         );
  CMX2X2 U3027 ( .A0(\memory[7][26] ), .A1(out_new[26]), .S(N3107), .Z(n1849)
         );
  CMX2X2 U3028 ( .A0(\memory[7][25] ), .A1(out_new[25]), .S(N3107), .Z(n1850)
         );
  CMX2X2 U3029 ( .A0(\memory[7][24] ), .A1(out_new[24]), .S(N3107), .Z(n1851)
         );
  CMX2X2 U3030 ( .A0(\memory[7][23] ), .A1(out_new[23]), .S(N3107), .Z(n1852)
         );
  CMX2X2 U3031 ( .A0(\memory[7][22] ), .A1(out_new[22]), .S(N3107), .Z(n1853)
         );
  CMX2X2 U3032 ( .A0(\memory[7][21] ), .A1(out_new[21]), .S(N3107), .Z(n1854)
         );
  CMX2X2 U3033 ( .A0(\memory[7][20] ), .A1(out_new[20]), .S(N3107), .Z(n1855)
         );
  CMX2X2 U3034 ( .A0(\memory[7][19] ), .A1(out_new[19]), .S(N3107), .Z(n1856)
         );
  CMX2X2 U3035 ( .A0(\memory[7][18] ), .A1(out_new[18]), .S(N3107), .Z(n1857)
         );
  CMX2X2 U3036 ( .A0(\memory[7][17] ), .A1(out_new[17]), .S(N3107), .Z(n1858)
         );
  CMX2X2 U3037 ( .A0(\memory[7][16] ), .A1(out_new[16]), .S(N3107), .Z(n1859)
         );
  CMX2X2 U3038 ( .A0(\memory[7][15] ), .A1(out_new[15]), .S(N3107), .Z(n1860)
         );
  CMX2X2 U3039 ( .A0(\memory[7][14] ), .A1(out_new[14]), .S(N3107), .Z(n1861)
         );
  CMX2X2 U3040 ( .A0(\memory[7][13] ), .A1(out_new[13]), .S(N3107), .Z(n1862)
         );
  CMX2X2 U3041 ( .A0(\memory[7][12] ), .A1(out_new[12]), .S(N3107), .Z(n1863)
         );
  CMX2X2 U3042 ( .A0(\memory[7][11] ), .A1(out_new[11]), .S(N3107), .Z(n1864)
         );
  CMX2X2 U3043 ( .A0(\memory[7][10] ), .A1(out_new[10]), .S(N3107), .Z(n1865)
         );
  CMX2X2 U3044 ( .A0(\memory[7][9] ), .A1(out_new[9]), .S(N3107), .Z(n1866) );
  CMX2X2 U3045 ( .A0(\memory[7][8] ), .A1(out_new[8]), .S(N3107), .Z(n1867) );
  CMX2X2 U3046 ( .A0(\memory[7][7] ), .A1(out_new[7]), .S(N3107), .Z(n1868) );
  CMX2X2 U3047 ( .A0(\memory[7][6] ), .A1(out_new[6]), .S(N3107), .Z(n1869) );
  CMX2X2 U3048 ( .A0(\memory[7][5] ), .A1(out_new[5]), .S(N3107), .Z(n1870) );
  CMX2X2 U3049 ( .A0(\memory[7][4] ), .A1(out_new[4]), .S(N3107), .Z(n1871) );
  CMX2X2 U3050 ( .A0(\memory[7][3] ), .A1(out_new[3]), .S(N3107), .Z(n1872) );
  CMX2X2 U3051 ( .A0(\memory[7][2] ), .A1(out_new[2]), .S(N3107), .Z(n1873) );
  CMX2X2 U3052 ( .A0(\memory[7][1] ), .A1(out_new[1]), .S(N3107), .Z(n1874) );
  CMX2X2 U3053 ( .A0(\memory[7][0] ), .A1(out_new[0]), .S(N3107), .Z(n1875) );
  CMX2X4 U3054 ( .A0(lenout[5]), .A1(N44), .S(N4960), .Z(n2452) );
  CMX2X4 U3055 ( .A0(lenout[6]), .A1(N43), .S(N4960), .Z(n2453) );
  CMX2X4 U3056 ( .A0(lenout[4]), .A1(N45), .S(N4960), .Z(n2451) );
  CMX2X4 U3057 ( .A0(lenout[3]), .A1(N46), .S(N4960), .Z(n2450) );
  CMX2X4 U3058 ( .A0(lenout[2]), .A1(N47), .S(N4960), .Z(n2449) );
  CMX2X4 U3059 ( .A0(lenout[1]), .A1(N48), .S(N4960), .Z(n2448) );
  CMX2X4 U3060 ( .A0(lenout[0]), .A1(N49), .S(N4960), .Z(n2447) );
  CMX2X4 U3061 ( .A0(dataout[63]), .A1(N50), .S(N4960), .Z(n2446) );
  CMX2X4 U3062 ( .A0(dataout[62]), .A1(N51), .S(N4960), .Z(n2445) );
  CMX2X4 U3063 ( .A0(dataout[61]), .A1(N52), .S(N4960), .Z(n2444) );
  CMX2X4 U3064 ( .A0(dataout[60]), .A1(N53), .S(N4960), .Z(n2443) );
  CMX2X4 U3065 ( .A0(dataout[59]), .A1(N54), .S(N4960), .Z(n2442) );
  CMX2X4 U3066 ( .A0(dataout[58]), .A1(N55), .S(N4960), .Z(n2441) );
  CMX2X4 U3067 ( .A0(dataout[57]), .A1(N56), .S(N4960), .Z(n2440) );
  CMX2X4 U3068 ( .A0(dataout[56]), .A1(N57), .S(N4960), .Z(n2439) );
  CMX2X4 U3069 ( .A0(dataout[55]), .A1(N58), .S(N4960), .Z(n2438) );
  CMX2X4 U3070 ( .A0(dataout[54]), .A1(N59), .S(N4960), .Z(n2437) );
  CMX2X4 U3071 ( .A0(dataout[53]), .A1(N60), .S(N4960), .Z(n2436) );
  CMX2X4 U3072 ( .A0(dataout[52]), .A1(N61), .S(N4960), .Z(n2435) );
  CMX2X4 U3073 ( .A0(dataout[51]), .A1(N62), .S(N4960), .Z(n2434) );
  CMX2X4 U3074 ( .A0(dataout[50]), .A1(N63), .S(N4960), .Z(n2433) );
  CMX2X4 U3075 ( .A0(dataout[49]), .A1(N64), .S(N4960), .Z(n2432) );
  CMX2X4 U3076 ( .A0(dataout[48]), .A1(N65), .S(N4960), .Z(n2431) );
  CMX2X4 U3077 ( .A0(dataout[47]), .A1(N66), .S(N4960), .Z(n2430) );
  CMX2X4 U3078 ( .A0(dataout[46]), .A1(N67), .S(N4960), .Z(n2429) );
  CMX2X4 U3079 ( .A0(dataout[45]), .A1(N68), .S(N4960), .Z(n2428) );
  CMX2X4 U3080 ( .A0(dataout[44]), .A1(N69), .S(N4960), .Z(n2427) );
  CMX2X4 U3081 ( .A0(dataout[43]), .A1(N70), .S(N4960), .Z(n2426) );
  CMX2X4 U3082 ( .A0(dataout[42]), .A1(N71), .S(N4960), .Z(n2425) );
  CMX2X4 U3083 ( .A0(dataout[41]), .A1(N72), .S(N4960), .Z(n2424) );
  CMX2X4 U3084 ( .A0(dataout[40]), .A1(N73), .S(N4960), .Z(n2423) );
  CMX2X4 U3085 ( .A0(dataout[39]), .A1(N74), .S(N4960), .Z(n2422) );
  CMX2X4 U3086 ( .A0(dataout[38]), .A1(N75), .S(N4960), .Z(n2421) );
  CMX2X4 U3087 ( .A0(dataout[37]), .A1(N76), .S(N4960), .Z(n2420) );
  CMX2X4 U3088 ( .A0(dataout[36]), .A1(N77), .S(N4960), .Z(n2419) );
  CMX2X4 U3089 ( .A0(dataout[35]), .A1(N78), .S(N4960), .Z(n2418) );
  CMX2X4 U3090 ( .A0(dataout[34]), .A1(N79), .S(N4960), .Z(n2417) );
  CMX2X4 U3091 ( .A0(dataout[33]), .A1(N80), .S(N4960), .Z(n2416) );
  CMX2X4 U3092 ( .A0(dataout[32]), .A1(N81), .S(N4960), .Z(n2415) );
  CMX2X4 U3093 ( .A0(dataout[31]), .A1(N82), .S(N4960), .Z(n2414) );
  CMX2X4 U3094 ( .A0(dataout[30]), .A1(N83), .S(N4960), .Z(n2413) );
  CMX2X4 U3095 ( .A0(dataout[29]), .A1(N84), .S(N4960), .Z(n2412) );
  CMX2X4 U3096 ( .A0(dataout[28]), .A1(N85), .S(N4960), .Z(n2411) );
  CMX2X4 U3097 ( .A0(dataout[27]), .A1(N86), .S(N4960), .Z(n2410) );
  CMX2X4 U3098 ( .A0(dataout[26]), .A1(N87), .S(N4960), .Z(n2409) );
  CMX2X4 U3099 ( .A0(dataout[25]), .A1(N88), .S(N4960), .Z(n2408) );
  CMX2X4 U3100 ( .A0(dataout[24]), .A1(N89), .S(N4960), .Z(n2407) );
  CMX2X4 U3101 ( .A0(dataout[23]), .A1(N90), .S(N4960), .Z(n2406) );
  CMX2X4 U3102 ( .A0(dataout[22]), .A1(N91), .S(N4960), .Z(n2405) );
  CMX2X4 U3103 ( .A0(dataout[21]), .A1(N92), .S(N4960), .Z(n2404) );
  CMX2X4 U3104 ( .A0(dataout[20]), .A1(N93), .S(N4960), .Z(n2403) );
  CMX2X4 U3105 ( .A0(dataout[19]), .A1(N94), .S(N4960), .Z(n2402) );
  CMX2X4 U3106 ( .A0(dataout[18]), .A1(N95), .S(N4960), .Z(n2401) );
  CMX2X4 U3107 ( .A0(dataout[17]), .A1(N96), .S(N4960), .Z(n2400) );
  CMX2X4 U3108 ( .A0(dataout[16]), .A1(N97), .S(N4960), .Z(n2399) );
  CMX2X4 U3109 ( .A0(dataout[15]), .A1(N98), .S(N4960), .Z(n2398) );
  CMX2X4 U3110 ( .A0(dataout[14]), .A1(N99), .S(N4960), .Z(n2397) );
  CMX2X4 U3111 ( .A0(dataout[13]), .A1(N100), .S(N4960), .Z(n2396) );
  CMX2X4 U3112 ( .A0(dataout[12]), .A1(N101), .S(N4960), .Z(n2395) );
  CMX2X4 U3113 ( .A0(dataout[11]), .A1(N102), .S(N4960), .Z(n2394) );
  CMX2X4 U3114 ( .A0(dataout[10]), .A1(N103), .S(N4960), .Z(n2393) );
  CMX2X4 U3115 ( .A0(dataout[9]), .A1(N104), .S(N4960), .Z(n2392) );
  CMX2X4 U3116 ( .A0(dataout[8]), .A1(N105), .S(N4960), .Z(n2391) );
  CMX2X4 U3117 ( .A0(dataout[7]), .A1(N106), .S(N4960), .Z(n2390) );
  CMX2X4 U3118 ( .A0(dataout[6]), .A1(N107), .S(N4960), .Z(n2389) );
  CMX2X4 U3119 ( .A0(dataout[5]), .A1(N108), .S(N4960), .Z(n2388) );
  CMX2X4 U3120 ( .A0(dataout[4]), .A1(N109), .S(N4960), .Z(n2387) );
  CMX2X4 U3121 ( .A0(dataout[3]), .A1(N110), .S(N4960), .Z(n2386) );
  CMX2X4 U3122 ( .A0(dataout[2]), .A1(N111), .S(N4960), .Z(n2385) );
  CMX2X4 U3123 ( .A0(dataout[1]), .A1(N112), .S(N4960), .Z(n2384) );
  CMX2X4 U3124 ( .A0(dataout[0]), .A1(N113), .S(N4960), .Z(n2383) );
  CMX2X2 U3125 ( .A0(\memory[27][62] ), .A1(out_new[62]), .S(N4527), .Z(n393)
         );
  CMX2X2 U3126 ( .A0(\memory[23][62] ), .A1(out_new[62]), .S(N4243), .Z(n677)
         );
  CMX2X2 U3127 ( .A0(\memory[19][62] ), .A1(out_new[62]), .S(N3959), .Z(n961)
         );
  CMX2X2 U3128 ( .A0(\memory[15][62] ), .A1(out_new[62]), .S(N3675), .Z(n1245)
         );
  CNIVXL U3129 ( .A(out[62]), .Z(n2536) );
  CNIVX1 U3130 ( .A(out[61]), .Z(n2537) );
  CNIVX1 U3131 ( .A(out[60]), .Z(n2538) );
  CNIVX1 U3132 ( .A(out[59]), .Z(n2539) );
  CNIVX1 U3133 ( .A(out[58]), .Z(n2540) );
  CNIVX1 U3134 ( .A(out[57]), .Z(n2541) );
  CNIVX1 U3135 ( .A(out[56]), .Z(n2542) );
  CNIVX1 U3136 ( .A(out[55]), .Z(n2543) );
  CNIVX1 U3137 ( .A(out[54]), .Z(n2544) );
  CNIVX1 U3138 ( .A(out[53]), .Z(n2545) );
  CNIVX1 U3139 ( .A(out[52]), .Z(n2546) );
  CNIVX1 U3140 ( .A(out[51]), .Z(n2547) );
  CNIVX1 U3141 ( .A(out[50]), .Z(n2548) );
  CNIVX1 U3142 ( .A(out[49]), .Z(n2549) );
  CNIVX1 U3143 ( .A(out[48]), .Z(n2550) );
  CNIVX1 U3144 ( .A(out[47]), .Z(n2551) );
  CNIVX1 U3145 ( .A(out[46]), .Z(n2552) );
  CNIVX1 U3146 ( .A(out[45]), .Z(n2553) );
  CNIVX1 U3147 ( .A(out[44]), .Z(n2554) );
  CNIVX1 U3148 ( .A(out[43]), .Z(n2555) );
  CNIVX1 U3149 ( .A(out[42]), .Z(n2556) );
  CNIVX1 U3150 ( .A(out[41]), .Z(n2557) );
  CNIVX1 U3151 ( .A(out[40]), .Z(n2558) );
  CNIVX1 U3152 ( .A(out[39]), .Z(n2559) );
  CNIVX1 U3153 ( .A(out[38]), .Z(n2560) );
  CNIVX1 U3154 ( .A(out[37]), .Z(n2561) );
  CNIVX1 U3155 ( .A(out[36]), .Z(n2562) );
  CNIVX1 U3156 ( .A(out[35]), .Z(n2563) );
  CNIVX1 U3157 ( .A(out[34]), .Z(n2564) );
  CNIVX1 U3158 ( .A(out[33]), .Z(n2565) );
  CNIVX1 U3159 ( .A(out[32]), .Z(n2566) );
  CNIVX1 U3160 ( .A(out[31]), .Z(n2567) );
  CNIVX1 U3161 ( .A(out[30]), .Z(n2568) );
  CNIVX1 U3162 ( .A(out[29]), .Z(n2569) );
  CNIVX1 U3163 ( .A(out[28]), .Z(n2570) );
  CNIVX1 U3164 ( .A(out[27]), .Z(n2571) );
  CNIVX1 U3165 ( .A(out[26]), .Z(n2572) );
  CNIVX1 U3166 ( .A(out[25]), .Z(n2573) );
  CNIVX1 U3167 ( .A(out[24]), .Z(n2574) );
  CNIVX1 U3168 ( .A(out[23]), .Z(n2575) );
  CNIVX1 U3169 ( .A(out[22]), .Z(n2576) );
  CNIVX1 U3170 ( .A(out[21]), .Z(n2577) );
  CNIVX1 U3171 ( .A(out[20]), .Z(n2578) );
  CNIVX1 U3172 ( .A(out[19]), .Z(n2579) );
  CNIVX1 U3173 ( .A(out[18]), .Z(n2580) );
  CNIVX1 U3174 ( .A(out[17]), .Z(n2581) );
  CNIVX1 U3175 ( .A(out[16]), .Z(n2582) );
  CNIVX1 U3176 ( .A(out[15]), .Z(n2583) );
  CNIVX1 U3177 ( .A(out[14]), .Z(n2584) );
  CNIVX1 U3178 ( .A(out[13]), .Z(n2585) );
  CNIVX1 U3179 ( .A(out[12]), .Z(n2586) );
  CNIVX1 U3180 ( .A(out[11]), .Z(n2587) );
  CNIVX1 U3181 ( .A(out[10]), .Z(n2588) );
  CNIVX1 U3182 ( .A(out[9]), .Z(n2589) );
  CNIVX1 U3183 ( .A(out[8]), .Z(n2590) );
  CNIVX1 U3184 ( .A(out[7]), .Z(n2591) );
  CNIVX1 U3185 ( .A(out[6]), .Z(n2592) );
  CNIVX1 U3186 ( .A(out[5]), .Z(n2593) );
  CNIVX1 U3187 ( .A(out[4]), .Z(n2594) );
  CNIVX1 U3188 ( .A(out[3]), .Z(n2595) );
  CNIVX1 U3189 ( .A(out[2]), .Z(n2596) );
  CNIVX1 U3190 ( .A(out[1]), .Z(n2597) );
  CNIVX1 U3191 ( .A(out[0]), .Z(n2598) );
  CNIVX1 U3192 ( .A(lout[0]), .Z(n2599) );
  CMX2X2 U3193 ( .A0(\memory[27][63] ), .A1(out_new[63]), .S(N4527), .Z(n392)
         );
  CMX2X2 U3194 ( .A0(\memory[27][61] ), .A1(out_new[61]), .S(N4527), .Z(n394)
         );
  CMX2X2 U3195 ( .A0(\memory[27][60] ), .A1(out_new[60]), .S(N4527), .Z(n395)
         );
  CMX2X2 U3196 ( .A0(\memory[27][59] ), .A1(out_new[59]), .S(N4527), .Z(n396)
         );
  CMX2X2 U3197 ( .A0(\memory[27][58] ), .A1(out_new[58]), .S(N4527), .Z(n397)
         );
  CMX2X2 U3198 ( .A0(\memory[27][57] ), .A1(out_new[57]), .S(N4527), .Z(n398)
         );
  CMX2X2 U3199 ( .A0(\memory[27][56] ), .A1(out_new[56]), .S(N4527), .Z(n399)
         );
  CMX2X2 U3200 ( .A0(\memory[27][55] ), .A1(out_new[55]), .S(N4527), .Z(n400)
         );
  CMX2X2 U3201 ( .A0(\memory[27][54] ), .A1(out_new[54]), .S(N4527), .Z(n401)
         );
  CMX2X2 U3202 ( .A0(\memory[27][53] ), .A1(out_new[53]), .S(N4527), .Z(n402)
         );
  CMX2X2 U3203 ( .A0(\memory[27][52] ), .A1(out_new[52]), .S(N4527), .Z(n403)
         );
  CMX2X2 U3204 ( .A0(\memory[27][51] ), .A1(out_new[51]), .S(N4527), .Z(n404)
         );
  CMX2X2 U3205 ( .A0(\memory[27][50] ), .A1(out_new[50]), .S(N4527), .Z(n405)
         );
  CMX2X2 U3206 ( .A0(\memory[27][49] ), .A1(out_new[49]), .S(N4527), .Z(n406)
         );
  CMX2X2 U3207 ( .A0(\memory[27][48] ), .A1(out_new[48]), .S(N4527), .Z(n407)
         );
  CMX2X2 U3208 ( .A0(\memory[27][47] ), .A1(out_new[47]), .S(N4527), .Z(n408)
         );
  CMX2X2 U3209 ( .A0(\memory[27][46] ), .A1(out_new[46]), .S(N4527), .Z(n409)
         );
  CMX2X2 U3210 ( .A0(\memory[27][45] ), .A1(out_new[45]), .S(N4527), .Z(n410)
         );
  CMX2X2 U3211 ( .A0(\memory[27][44] ), .A1(out_new[44]), .S(N4527), .Z(n411)
         );
  CMX2X2 U3212 ( .A0(\memory[27][43] ), .A1(out_new[43]), .S(N4527), .Z(n412)
         );
  CMX2X2 U3213 ( .A0(\memory[27][42] ), .A1(out_new[42]), .S(N4527), .Z(n413)
         );
  CMX2X2 U3214 ( .A0(\memory[27][41] ), .A1(out_new[41]), .S(N4527), .Z(n414)
         );
  CMX2X2 U3215 ( .A0(\memory[27][40] ), .A1(out_new[40]), .S(N4527), .Z(n415)
         );
  CMX2X2 U3216 ( .A0(\memory[27][39] ), .A1(out_new[39]), .S(N4527), .Z(n416)
         );
  CMX2X2 U3217 ( .A0(\memory[27][38] ), .A1(out_new[38]), .S(N4527), .Z(n417)
         );
  CMX2X2 U3218 ( .A0(\memory[27][37] ), .A1(out_new[37]), .S(N4527), .Z(n418)
         );
  CMX2X2 U3219 ( .A0(\memory[27][36] ), .A1(out_new[36]), .S(N4527), .Z(n419)
         );
  CMX2X2 U3220 ( .A0(\memory[27][35] ), .A1(out_new[35]), .S(N4527), .Z(n420)
         );
  CMX2X2 U3221 ( .A0(\memory[27][34] ), .A1(out_new[34]), .S(N4527), .Z(n421)
         );
  CMX2X2 U3222 ( .A0(\memory[27][33] ), .A1(out_new[33]), .S(N4527), .Z(n422)
         );
  CMX2X2 U3223 ( .A0(\memory[27][32] ), .A1(out_new[32]), .S(N4527), .Z(n423)
         );
  CMX2X2 U3224 ( .A0(\memory[27][31] ), .A1(out_new[31]), .S(N4527), .Z(n424)
         );
  CMX2X2 U3225 ( .A0(\memory[27][30] ), .A1(out_new[30]), .S(N4527), .Z(n425)
         );
  CMX2X2 U3226 ( .A0(\memory[27][29] ), .A1(out_new[29]), .S(N4527), .Z(n426)
         );
  CMX2X2 U3227 ( .A0(\memory[27][28] ), .A1(out_new[28]), .S(N4527), .Z(n427)
         );
  CMX2X2 U3228 ( .A0(\memory[27][27] ), .A1(out_new[27]), .S(N4527), .Z(n428)
         );
  CMX2X2 U3229 ( .A0(\memory[27][26] ), .A1(out_new[26]), .S(N4527), .Z(n429)
         );
  CMX2X2 U3230 ( .A0(\memory[27][25] ), .A1(out_new[25]), .S(N4527), .Z(n430)
         );
  CMX2X2 U3231 ( .A0(\memory[27][24] ), .A1(out_new[24]), .S(N4527), .Z(n431)
         );
  CMX2X2 U3232 ( .A0(\memory[27][23] ), .A1(out_new[23]), .S(N4527), .Z(n432)
         );
  CMX2X2 U3233 ( .A0(\memory[27][22] ), .A1(out_new[22]), .S(N4527), .Z(n433)
         );
  CMX2X2 U3234 ( .A0(\memory[27][21] ), .A1(out_new[21]), .S(N4527), .Z(n434)
         );
  CMX2X2 U3235 ( .A0(\memory[27][20] ), .A1(out_new[20]), .S(N4527), .Z(n435)
         );
  CMX2X2 U3236 ( .A0(\memory[27][19] ), .A1(out_new[19]), .S(N4527), .Z(n436)
         );
  CMX2X2 U3237 ( .A0(\memory[27][18] ), .A1(out_new[18]), .S(N4527), .Z(n437)
         );
  CMX2X2 U3238 ( .A0(\memory[27][17] ), .A1(out_new[17]), .S(N4527), .Z(n438)
         );
  CMX2X2 U3239 ( .A0(\memory[27][16] ), .A1(out_new[16]), .S(N4527), .Z(n439)
         );
  CMX2X2 U3240 ( .A0(\memory[27][15] ), .A1(out_new[15]), .S(N4527), .Z(n440)
         );
  CMX2X2 U3241 ( .A0(\memory[27][14] ), .A1(out_new[14]), .S(N4527), .Z(n441)
         );
  CMX2X2 U3242 ( .A0(\memory[27][13] ), .A1(out_new[13]), .S(N4527), .Z(n442)
         );
  CMX2X2 U3243 ( .A0(\memory[27][12] ), .A1(out_new[12]), .S(N4527), .Z(n443)
         );
  CMX2X2 U3244 ( .A0(\memory[27][11] ), .A1(out_new[11]), .S(N4527), .Z(n444)
         );
  CMX2X2 U3245 ( .A0(\memory[27][10] ), .A1(out_new[10]), .S(N4527), .Z(n445)
         );
  CMX2X2 U3246 ( .A0(\memory[27][9] ), .A1(out_new[9]), .S(N4527), .Z(n446) );
  CMX2X2 U3247 ( .A0(\memory[27][8] ), .A1(out_new[8]), .S(N4527), .Z(n447) );
  CMX2X2 U3248 ( .A0(\memory[27][7] ), .A1(out_new[7]), .S(N4527), .Z(n448) );
  CMX2X2 U3249 ( .A0(\memory[27][6] ), .A1(out_new[6]), .S(N4527), .Z(n449) );
  CMX2X2 U3250 ( .A0(\memory[27][5] ), .A1(out_new[5]), .S(N4527), .Z(n450) );
  CMX2X2 U3251 ( .A0(\memory[27][4] ), .A1(out_new[4]), .S(N4527), .Z(n451) );
  CMX2X2 U3252 ( .A0(\memory[27][3] ), .A1(out_new[3]), .S(N4527), .Z(n452) );
  CMX2X2 U3253 ( .A0(\memory[27][2] ), .A1(out_new[2]), .S(N4527), .Z(n453) );
  CMX2X2 U3254 ( .A0(\memory[27][1] ), .A1(out_new[1]), .S(N4527), .Z(n454) );
  CMX2X2 U3255 ( .A0(\memory[27][0] ), .A1(out_new[0]), .S(N4527), .Z(n455) );
  CMX2X2 U3256 ( .A0(\memory[23][63] ), .A1(out_new[63]), .S(N4243), .Z(n676)
         );
  CMX2X2 U3257 ( .A0(\memory[23][61] ), .A1(out_new[61]), .S(N4243), .Z(n678)
         );
  CMX2X2 U3258 ( .A0(\memory[23][60] ), .A1(out_new[60]), .S(N4243), .Z(n679)
         );
  CMX2X2 U3259 ( .A0(\memory[23][59] ), .A1(out_new[59]), .S(N4243), .Z(n680)
         );
  CMX2X2 U3260 ( .A0(\memory[23][58] ), .A1(out_new[58]), .S(N4243), .Z(n681)
         );
  CMX2X2 U3261 ( .A0(\memory[23][57] ), .A1(out_new[57]), .S(N4243), .Z(n682)
         );
  CMX2X2 U3262 ( .A0(\memory[23][56] ), .A1(out_new[56]), .S(N4243), .Z(n683)
         );
  CMX2X2 U3263 ( .A0(\memory[23][55] ), .A1(out_new[55]), .S(N4243), .Z(n684)
         );
  CMX2X2 U3264 ( .A0(\memory[23][54] ), .A1(out_new[54]), .S(N4243), .Z(n685)
         );
  CMX2X2 U3265 ( .A0(\memory[23][53] ), .A1(out_new[53]), .S(N4243), .Z(n686)
         );
  CMX2X2 U3266 ( .A0(\memory[23][52] ), .A1(out_new[52]), .S(N4243), .Z(n687)
         );
  CMX2X2 U3267 ( .A0(\memory[23][51] ), .A1(out_new[51]), .S(N4243), .Z(n688)
         );
  CMX2X2 U3268 ( .A0(\memory[23][50] ), .A1(out_new[50]), .S(N4243), .Z(n689)
         );
  CMX2X2 U3269 ( .A0(\memory[23][49] ), .A1(out_new[49]), .S(N4243), .Z(n690)
         );
  CMX2X2 U3270 ( .A0(\memory[23][48] ), .A1(out_new[48]), .S(N4243), .Z(n691)
         );
  CMX2X2 U3271 ( .A0(\memory[23][47] ), .A1(out_new[47]), .S(N4243), .Z(n692)
         );
  CMX2X2 U3272 ( .A0(\memory[23][46] ), .A1(out_new[46]), .S(N4243), .Z(n693)
         );
  CMX2X2 U3273 ( .A0(\memory[23][45] ), .A1(out_new[45]), .S(N4243), .Z(n694)
         );
  CMX2X2 U3274 ( .A0(\memory[23][44] ), .A1(out_new[44]), .S(N4243), .Z(n695)
         );
  CMX2X2 U3275 ( .A0(\memory[23][43] ), .A1(out_new[43]), .S(N4243), .Z(n696)
         );
  CMX2X2 U3276 ( .A0(\memory[23][42] ), .A1(out_new[42]), .S(N4243), .Z(n697)
         );
  CMX2X2 U3277 ( .A0(\memory[23][41] ), .A1(out_new[41]), .S(N4243), .Z(n698)
         );
  CMX2X2 U3278 ( .A0(\memory[23][40] ), .A1(out_new[40]), .S(N4243), .Z(n699)
         );
  CMX2X2 U3279 ( .A0(\memory[23][39] ), .A1(out_new[39]), .S(N4243), .Z(n700)
         );
  CMX2X2 U3280 ( .A0(\memory[23][38] ), .A1(out_new[38]), .S(N4243), .Z(n701)
         );
  CMX2X2 U3281 ( .A0(\memory[23][37] ), .A1(out_new[37]), .S(N4243), .Z(n702)
         );
  CMX2X2 U3282 ( .A0(\memory[23][36] ), .A1(out_new[36]), .S(N4243), .Z(n703)
         );
  CMX2X2 U3283 ( .A0(\memory[23][35] ), .A1(out_new[35]), .S(N4243), .Z(n704)
         );
  CMX2X2 U3284 ( .A0(\memory[23][34] ), .A1(out_new[34]), .S(N4243), .Z(n705)
         );
  CMX2X2 U3285 ( .A0(\memory[23][33] ), .A1(out_new[33]), .S(N4243), .Z(n706)
         );
  CMX2X2 U3286 ( .A0(\memory[23][32] ), .A1(out_new[32]), .S(N4243), .Z(n707)
         );
  CMX2X2 U3287 ( .A0(\memory[23][31] ), .A1(out_new[31]), .S(N4243), .Z(n708)
         );
  CMX2X2 U3288 ( .A0(\memory[23][30] ), .A1(out_new[30]), .S(N4243), .Z(n709)
         );
  CMX2X2 U3289 ( .A0(\memory[23][29] ), .A1(out_new[29]), .S(N4243), .Z(n710)
         );
  CMX2X2 U3290 ( .A0(\memory[23][28] ), .A1(out_new[28]), .S(N4243), .Z(n711)
         );
  CMX2X2 U3291 ( .A0(\memory[23][27] ), .A1(out_new[27]), .S(N4243), .Z(n712)
         );
  CMX2X2 U3292 ( .A0(\memory[23][26] ), .A1(out_new[26]), .S(N4243), .Z(n713)
         );
  CMX2X2 U3293 ( .A0(\memory[23][25] ), .A1(out_new[25]), .S(N4243), .Z(n714)
         );
  CMX2X2 U3294 ( .A0(\memory[23][24] ), .A1(out_new[24]), .S(N4243), .Z(n715)
         );
  CMX2X2 U3295 ( .A0(\memory[23][23] ), .A1(out_new[23]), .S(N4243), .Z(n716)
         );
  CMX2X2 U3296 ( .A0(\memory[23][22] ), .A1(out_new[22]), .S(N4243), .Z(n717)
         );
  CMX2X2 U3297 ( .A0(\memory[23][21] ), .A1(out_new[21]), .S(N4243), .Z(n718)
         );
  CMX2X2 U3298 ( .A0(\memory[23][20] ), .A1(out_new[20]), .S(N4243), .Z(n719)
         );
  CMX2X2 U3299 ( .A0(\memory[23][19] ), .A1(out_new[19]), .S(N4243), .Z(n720)
         );
  CMX2X2 U3300 ( .A0(\memory[23][18] ), .A1(out_new[18]), .S(N4243), .Z(n721)
         );
  CMX2X2 U3301 ( .A0(\memory[23][17] ), .A1(out_new[17]), .S(N4243), .Z(n722)
         );
  CMX2X2 U3302 ( .A0(\memory[23][16] ), .A1(out_new[16]), .S(N4243), .Z(n723)
         );
  CMX2X2 U3303 ( .A0(\memory[23][15] ), .A1(out_new[15]), .S(N4243), .Z(n724)
         );
  CMX2X2 U3304 ( .A0(\memory[23][14] ), .A1(out_new[14]), .S(N4243), .Z(n725)
         );
  CMX2X2 U3305 ( .A0(\memory[23][13] ), .A1(out_new[13]), .S(N4243), .Z(n726)
         );
  CMX2X2 U3306 ( .A0(\memory[23][12] ), .A1(out_new[12]), .S(N4243), .Z(n727)
         );
  CMX2X2 U3307 ( .A0(\memory[23][11] ), .A1(out_new[11]), .S(N4243), .Z(n728)
         );
  CMX2X2 U3308 ( .A0(\memory[23][10] ), .A1(out_new[10]), .S(N4243), .Z(n729)
         );
  CMX2X2 U3309 ( .A0(\memory[23][9] ), .A1(out_new[9]), .S(N4243), .Z(n730) );
  CMX2X2 U3310 ( .A0(\memory[23][8] ), .A1(out_new[8]), .S(N4243), .Z(n731) );
  CMX2X2 U3311 ( .A0(\memory[23][7] ), .A1(out_new[7]), .S(N4243), .Z(n732) );
  CMX2X2 U3312 ( .A0(\memory[23][6] ), .A1(out_new[6]), .S(N4243), .Z(n733) );
  CMX2X2 U3313 ( .A0(\memory[23][5] ), .A1(out_new[5]), .S(N4243), .Z(n734) );
  CMX2X2 U3314 ( .A0(\memory[23][4] ), .A1(out_new[4]), .S(N4243), .Z(n735) );
  CMX2X2 U3315 ( .A0(\memory[23][3] ), .A1(out_new[3]), .S(N4243), .Z(n736) );
  CMX2X2 U3316 ( .A0(\memory[23][2] ), .A1(out_new[2]), .S(N4243), .Z(n737) );
  CMX2X2 U3317 ( .A0(\memory[23][1] ), .A1(out_new[1]), .S(N4243), .Z(n738) );
  CMX2X2 U3318 ( .A0(\memory[23][0] ), .A1(out_new[0]), .S(N4243), .Z(n739) );
  CMX2X2 U3319 ( .A0(\memory[19][63] ), .A1(out_new[63]), .S(N3959), .Z(n960)
         );
  CMX2X2 U3320 ( .A0(\memory[19][61] ), .A1(out_new[61]), .S(N3959), .Z(n962)
         );
  CMX2X2 U3321 ( .A0(\memory[19][60] ), .A1(out_new[60]), .S(N3959), .Z(n963)
         );
  CMX2X2 U3322 ( .A0(\memory[19][59] ), .A1(out_new[59]), .S(N3959), .Z(n964)
         );
  CMX2X2 U3323 ( .A0(\memory[19][58] ), .A1(out_new[58]), .S(N3959), .Z(n965)
         );
  CMX2X2 U3324 ( .A0(\memory[19][57] ), .A1(out_new[57]), .S(N3959), .Z(n966)
         );
  CMX2X2 U3325 ( .A0(\memory[19][56] ), .A1(out_new[56]), .S(N3959), .Z(n967)
         );
  CMX2X2 U3326 ( .A0(\memory[19][55] ), .A1(out_new[55]), .S(N3959), .Z(n968)
         );
  CMX2X2 U3327 ( .A0(\memory[19][54] ), .A1(out_new[54]), .S(N3959), .Z(n969)
         );
  CMX2X2 U3328 ( .A0(\memory[19][53] ), .A1(out_new[53]), .S(N3959), .Z(n970)
         );
  CMX2X2 U3329 ( .A0(\memory[19][52] ), .A1(out_new[52]), .S(N3959), .Z(n971)
         );
  CMX2X2 U3330 ( .A0(\memory[19][51] ), .A1(out_new[51]), .S(N3959), .Z(n972)
         );
  CMX2X2 U3331 ( .A0(\memory[19][50] ), .A1(out_new[50]), .S(N3959), .Z(n973)
         );
  CMX2X2 U3332 ( .A0(\memory[19][49] ), .A1(out_new[49]), .S(N3959), .Z(n974)
         );
  CMX2X2 U3333 ( .A0(\memory[19][48] ), .A1(out_new[48]), .S(N3959), .Z(n975)
         );
  CMX2X2 U3334 ( .A0(\memory[19][47] ), .A1(out_new[47]), .S(N3959), .Z(n976)
         );
  CMX2X2 U3335 ( .A0(\memory[19][46] ), .A1(out_new[46]), .S(N3959), .Z(n977)
         );
  CMX2X2 U3336 ( .A0(\memory[19][45] ), .A1(out_new[45]), .S(N3959), .Z(n978)
         );
  CMX2X2 U3337 ( .A0(\memory[19][44] ), .A1(out_new[44]), .S(N3959), .Z(n979)
         );
  CMX2X2 U3338 ( .A0(\memory[19][43] ), .A1(out_new[43]), .S(N3959), .Z(n980)
         );
  CMX2X2 U3339 ( .A0(\memory[19][42] ), .A1(out_new[42]), .S(N3959), .Z(n981)
         );
  CMX2X2 U3340 ( .A0(\memory[19][41] ), .A1(out_new[41]), .S(N3959), .Z(n982)
         );
  CMX2X2 U3341 ( .A0(\memory[19][40] ), .A1(out_new[40]), .S(N3959), .Z(n983)
         );
  CMX2X2 U3342 ( .A0(\memory[19][39] ), .A1(out_new[39]), .S(N3959), .Z(n984)
         );
  CMX2X2 U3343 ( .A0(\memory[19][38] ), .A1(out_new[38]), .S(N3959), .Z(n985)
         );
  CMX2X2 U3344 ( .A0(\memory[19][37] ), .A1(out_new[37]), .S(N3959), .Z(n986)
         );
  CMX2X2 U3345 ( .A0(\memory[19][36] ), .A1(out_new[36]), .S(N3959), .Z(n987)
         );
  CMX2X2 U3346 ( .A0(\memory[19][35] ), .A1(out_new[35]), .S(N3959), .Z(n988)
         );
  CMX2X2 U3347 ( .A0(\memory[19][34] ), .A1(out_new[34]), .S(N3959), .Z(n989)
         );
  CMX2X2 U3348 ( .A0(\memory[19][33] ), .A1(out_new[33]), .S(N3959), .Z(n990)
         );
  CMX2X2 U3349 ( .A0(\memory[19][32] ), .A1(out_new[32]), .S(N3959), .Z(n991)
         );
  CMX2X2 U3350 ( .A0(\memory[19][31] ), .A1(out_new[31]), .S(N3959), .Z(n992)
         );
  CMX2X2 U3351 ( .A0(\memory[19][30] ), .A1(out_new[30]), .S(N3959), .Z(n993)
         );
  CMX2X2 U3352 ( .A0(\memory[19][29] ), .A1(out_new[29]), .S(N3959), .Z(n994)
         );
  CMX2X2 U3353 ( .A0(\memory[19][28] ), .A1(out_new[28]), .S(N3959), .Z(n995)
         );
  CMX2X2 U3354 ( .A0(\memory[19][27] ), .A1(out_new[27]), .S(N3959), .Z(n996)
         );
  CMX2X2 U3355 ( .A0(\memory[19][26] ), .A1(out_new[26]), .S(N3959), .Z(n997)
         );
  CMX2X2 U3356 ( .A0(\memory[19][25] ), .A1(out_new[25]), .S(N3959), .Z(n998)
         );
  CMX2X2 U3357 ( .A0(\memory[19][24] ), .A1(out_new[24]), .S(N3959), .Z(n999)
         );
  CMX2X2 U3358 ( .A0(\memory[19][23] ), .A1(out_new[23]), .S(N3959), .Z(n1000)
         );
  CMX2X2 U3359 ( .A0(\memory[19][22] ), .A1(out_new[22]), .S(N3959), .Z(n1001)
         );
  CMX2X2 U3360 ( .A0(\memory[19][21] ), .A1(out_new[21]), .S(N3959), .Z(n1002)
         );
  CMX2X2 U3361 ( .A0(\memory[19][20] ), .A1(out_new[20]), .S(N3959), .Z(n1003)
         );
  CMX2X2 U3362 ( .A0(\memory[19][19] ), .A1(out_new[19]), .S(N3959), .Z(n1004)
         );
  CMX2X2 U3363 ( .A0(\memory[19][18] ), .A1(out_new[18]), .S(N3959), .Z(n1005)
         );
  CMX2X2 U3364 ( .A0(\memory[19][17] ), .A1(out_new[17]), .S(N3959), .Z(n1006)
         );
  CMX2X2 U3365 ( .A0(\memory[19][16] ), .A1(out_new[16]), .S(N3959), .Z(n1007)
         );
  CMX2X2 U3366 ( .A0(\memory[19][15] ), .A1(out_new[15]), .S(N3959), .Z(n1008)
         );
  CMX2X2 U3367 ( .A0(\memory[19][14] ), .A1(out_new[14]), .S(N3959), .Z(n1009)
         );
  CMX2X2 U3368 ( .A0(\memory[19][13] ), .A1(out_new[13]), .S(N3959), .Z(n1010)
         );
  CMX2X2 U3369 ( .A0(\memory[19][12] ), .A1(out_new[12]), .S(N3959), .Z(n1011)
         );
  CMX2X2 U3370 ( .A0(\memory[19][11] ), .A1(out_new[11]), .S(N3959), .Z(n1012)
         );
  CMX2X2 U3371 ( .A0(\memory[19][10] ), .A1(out_new[10]), .S(N3959), .Z(n1013)
         );
  CMX2X2 U3372 ( .A0(\memory[19][9] ), .A1(out_new[9]), .S(N3959), .Z(n1014)
         );
  CMX2X2 U3373 ( .A0(\memory[19][8] ), .A1(out_new[8]), .S(N3959), .Z(n1015)
         );
  CMX2X2 U3374 ( .A0(\memory[19][7] ), .A1(out_new[7]), .S(N3959), .Z(n1016)
         );
  CMX2X2 U3375 ( .A0(\memory[19][6] ), .A1(out_new[6]), .S(N3959), .Z(n1017)
         );
  CMX2X2 U3376 ( .A0(\memory[19][5] ), .A1(out_new[5]), .S(N3959), .Z(n1018)
         );
  CMX2X2 U3377 ( .A0(\memory[19][4] ), .A1(out_new[4]), .S(N3959), .Z(n1019)
         );
  CMX2X2 U3378 ( .A0(\memory[19][3] ), .A1(out_new[3]), .S(N3959), .Z(n1020)
         );
  CMX2X2 U3379 ( .A0(\memory[19][2] ), .A1(out_new[2]), .S(N3959), .Z(n1021)
         );
  CMX2X2 U3380 ( .A0(\memory[19][1] ), .A1(out_new[1]), .S(N3959), .Z(n1022)
         );
  CMX2X2 U3381 ( .A0(\memory[19][0] ), .A1(out_new[0]), .S(N3959), .Z(n1023)
         );
  CMX2X2 U3382 ( .A0(\memory[15][63] ), .A1(out_new[63]), .S(N3675), .Z(n1244)
         );
  CMX2X2 U3383 ( .A0(\memory[15][61] ), .A1(out_new[61]), .S(N3675), .Z(n1246)
         );
  CMX2X2 U3384 ( .A0(\memory[15][60] ), .A1(out_new[60]), .S(N3675), .Z(n1247)
         );
  CMX2X2 U3385 ( .A0(\memory[15][59] ), .A1(out_new[59]), .S(N3675), .Z(n1248)
         );
  CMX2X2 U3386 ( .A0(\memory[15][58] ), .A1(out_new[58]), .S(N3675), .Z(n1249)
         );
  CMX2X2 U3387 ( .A0(\memory[15][57] ), .A1(out_new[57]), .S(N3675), .Z(n1250)
         );
  CMX2X2 U3388 ( .A0(\memory[15][56] ), .A1(out_new[56]), .S(N3675), .Z(n1251)
         );
  CMX2X2 U3389 ( .A0(\memory[15][55] ), .A1(out_new[55]), .S(N3675), .Z(n1252)
         );
  CMX2X2 U3390 ( .A0(\memory[15][54] ), .A1(out_new[54]), .S(N3675), .Z(n1253)
         );
  CMX2X2 U3391 ( .A0(\memory[15][53] ), .A1(out_new[53]), .S(N3675), .Z(n1254)
         );
  CMX2X2 U3392 ( .A0(\memory[15][52] ), .A1(out_new[52]), .S(N3675), .Z(n1255)
         );
  CMX2X2 U3393 ( .A0(\memory[15][51] ), .A1(out_new[51]), .S(N3675), .Z(n1256)
         );
  CMX2X2 U3394 ( .A0(\memory[15][50] ), .A1(out_new[50]), .S(N3675), .Z(n1257)
         );
  CMX2X2 U3395 ( .A0(\memory[15][49] ), .A1(out_new[49]), .S(N3675), .Z(n1258)
         );
  CMX2X2 U3396 ( .A0(\memory[15][48] ), .A1(out_new[48]), .S(N3675), .Z(n1259)
         );
  CMX2X2 U3397 ( .A0(\memory[15][47] ), .A1(out_new[47]), .S(N3675), .Z(n1260)
         );
  CMX2X2 U3398 ( .A0(\memory[15][46] ), .A1(out_new[46]), .S(N3675), .Z(n1261)
         );
  CMX2X2 U3399 ( .A0(\memory[15][45] ), .A1(out_new[45]), .S(N3675), .Z(n1262)
         );
  CMX2X2 U3400 ( .A0(\memory[15][44] ), .A1(out_new[44]), .S(N3675), .Z(n1263)
         );
  CMX2X2 U3401 ( .A0(\memory[15][43] ), .A1(out_new[43]), .S(N3675), .Z(n1264)
         );
  CMX2X2 U3402 ( .A0(\memory[15][42] ), .A1(out_new[42]), .S(N3675), .Z(n1265)
         );
  CMX2X2 U3403 ( .A0(\memory[15][41] ), .A1(out_new[41]), .S(N3675), .Z(n1266)
         );
  CMX2X2 U3404 ( .A0(\memory[15][40] ), .A1(out_new[40]), .S(N3675), .Z(n1267)
         );
  CMX2X2 U3405 ( .A0(\memory[15][39] ), .A1(out_new[39]), .S(N3675), .Z(n1268)
         );
  CMX2X2 U3406 ( .A0(\memory[15][38] ), .A1(out_new[38]), .S(N3675), .Z(n1269)
         );
  CMX2X2 U3407 ( .A0(\memory[15][37] ), .A1(out_new[37]), .S(N3675), .Z(n1270)
         );
  CMX2X2 U3408 ( .A0(\memory[15][36] ), .A1(out_new[36]), .S(N3675), .Z(n1271)
         );
  CMX2X2 U3409 ( .A0(\memory[15][35] ), .A1(out_new[35]), .S(N3675), .Z(n1272)
         );
  CMX2X2 U3410 ( .A0(\memory[15][34] ), .A1(out_new[34]), .S(N3675), .Z(n1273)
         );
  CMX2X2 U3411 ( .A0(\memory[15][33] ), .A1(out_new[33]), .S(N3675), .Z(n1274)
         );
  CMX2X2 U3412 ( .A0(\memory[15][32] ), .A1(out_new[32]), .S(N3675), .Z(n1275)
         );
  CMX2X2 U3413 ( .A0(\memory[15][31] ), .A1(out_new[31]), .S(N3675), .Z(n1276)
         );
  CMX2X2 U3414 ( .A0(\memory[15][30] ), .A1(out_new[30]), .S(N3675), .Z(n1277)
         );
  CMX2X2 U3415 ( .A0(\memory[15][29] ), .A1(out_new[29]), .S(N3675), .Z(n1278)
         );
  CMX2X2 U3416 ( .A0(\memory[15][28] ), .A1(out_new[28]), .S(N3675), .Z(n1279)
         );
  CMX2X2 U3417 ( .A0(\memory[15][27] ), .A1(out_new[27]), .S(N3675), .Z(n1280)
         );
  CMX2X2 U3418 ( .A0(\memory[15][26] ), .A1(out_new[26]), .S(N3675), .Z(n1281)
         );
  CMX2X2 U3419 ( .A0(\memory[15][25] ), .A1(out_new[25]), .S(N3675), .Z(n1282)
         );
  CMX2X2 U3420 ( .A0(\memory[15][24] ), .A1(out_new[24]), .S(N3675), .Z(n1283)
         );
  CMX2X2 U3421 ( .A0(\memory[15][23] ), .A1(out_new[23]), .S(N3675), .Z(n1284)
         );
  CMX2X2 U3422 ( .A0(\memory[15][22] ), .A1(out_new[22]), .S(N3675), .Z(n1285)
         );
  CMX2X2 U3423 ( .A0(\memory[15][21] ), .A1(out_new[21]), .S(N3675), .Z(n1286)
         );
  CMX2X2 U3424 ( .A0(\memory[15][20] ), .A1(out_new[20]), .S(N3675), .Z(n1287)
         );
  CMX2X2 U3425 ( .A0(\memory[15][19] ), .A1(out_new[19]), .S(N3675), .Z(n1288)
         );
  CMX2X2 U3426 ( .A0(\memory[15][18] ), .A1(out_new[18]), .S(N3675), .Z(n1289)
         );
  CMX2X2 U3427 ( .A0(\memory[15][17] ), .A1(out_new[17]), .S(N3675), .Z(n1290)
         );
  CMX2X2 U3428 ( .A0(\memory[15][16] ), .A1(out_new[16]), .S(N3675), .Z(n1291)
         );
  CMX2X2 U3429 ( .A0(\memory[15][15] ), .A1(out_new[15]), .S(N3675), .Z(n1292)
         );
  CMX2X2 U3430 ( .A0(\memory[15][14] ), .A1(out_new[14]), .S(N3675), .Z(n1293)
         );
  CMX2X2 U3431 ( .A0(\memory[15][13] ), .A1(out_new[13]), .S(N3675), .Z(n1294)
         );
  CMX2X2 U3432 ( .A0(\memory[15][12] ), .A1(out_new[12]), .S(N3675), .Z(n1295)
         );
  CMX2X2 U3433 ( .A0(\memory[15][11] ), .A1(out_new[11]), .S(N3675), .Z(n1296)
         );
  CMX2X2 U3434 ( .A0(\memory[15][10] ), .A1(out_new[10]), .S(N3675), .Z(n1297)
         );
  CMX2X2 U3435 ( .A0(\memory[15][9] ), .A1(out_new[9]), .S(N3675), .Z(n1298)
         );
  CMX2X2 U3436 ( .A0(\memory[15][8] ), .A1(out_new[8]), .S(N3675), .Z(n1299)
         );
  CMX2X2 U3437 ( .A0(\memory[15][7] ), .A1(out_new[7]), .S(N3675), .Z(n1300)
         );
  CMX2X2 U3438 ( .A0(\memory[15][6] ), .A1(out_new[6]), .S(N3675), .Z(n1301)
         );
  CMX2X2 U3439 ( .A0(\memory[15][5] ), .A1(out_new[5]), .S(N3675), .Z(n1302)
         );
  CMX2X2 U3440 ( .A0(\memory[15][4] ), .A1(out_new[4]), .S(N3675), .Z(n1303)
         );
  CMX2X2 U3441 ( .A0(\memory[15][3] ), .A1(out_new[3]), .S(N3675), .Z(n1304)
         );
  CMX2X2 U3442 ( .A0(\memory[15][2] ), .A1(out_new[2]), .S(N3675), .Z(n1305)
         );
  CMX2X2 U3443 ( .A0(\memory[15][1] ), .A1(out_new[1]), .S(N3675), .Z(n1306)
         );
  CMX2X2 U3444 ( .A0(\memory[15][0] ), .A1(out_new[0]), .S(N3675), .Z(n1307)
         );
  CMX2X2 U3445 ( .A0(\memory[30][63] ), .A1(out_new[63]), .S(N4740), .Z(n179)
         );
  CMX2X2 U3446 ( .A0(\memory[30][62] ), .A1(out_new[62]), .S(N4740), .Z(n180)
         );
  CMX2X2 U3447 ( .A0(\memory[30][61] ), .A1(out_new[61]), .S(N4740), .Z(n181)
         );
  CMX2X2 U3448 ( .A0(\memory[30][60] ), .A1(out_new[60]), .S(N4740), .Z(n182)
         );
  CMX2X2 U3449 ( .A0(\memory[30][59] ), .A1(out_new[59]), .S(N4740), .Z(n183)
         );
  CMX2X2 U3450 ( .A0(\memory[30][58] ), .A1(out_new[58]), .S(N4740), .Z(n184)
         );
  CMX2X2 U3451 ( .A0(\memory[30][57] ), .A1(out_new[57]), .S(N4740), .Z(n185)
         );
  CMX2X2 U3452 ( .A0(\memory[30][56] ), .A1(out_new[56]), .S(N4740), .Z(n186)
         );
  CMX2X2 U3453 ( .A0(\memory[30][55] ), .A1(out_new[55]), .S(N4740), .Z(n187)
         );
  CMX2X2 U3454 ( .A0(\memory[30][54] ), .A1(out_new[54]), .S(N4740), .Z(n188)
         );
  CMX2X2 U3455 ( .A0(\memory[30][53] ), .A1(out_new[53]), .S(N4740), .Z(n189)
         );
  CMX2X2 U3456 ( .A0(\memory[30][52] ), .A1(out_new[52]), .S(N4740), .Z(n190)
         );
  CMX2X2 U3457 ( .A0(\memory[30][51] ), .A1(out_new[51]), .S(N4740), .Z(n191)
         );
  CMX2X2 U3458 ( .A0(\memory[30][50] ), .A1(out_new[50]), .S(N4740), .Z(n192)
         );
  CMX2X2 U3459 ( .A0(\memory[30][49] ), .A1(out_new[49]), .S(N4740), .Z(n193)
         );
  CMX2X2 U3460 ( .A0(\memory[30][48] ), .A1(out_new[48]), .S(N4740), .Z(n194)
         );
  CMX2X2 U3461 ( .A0(\memory[30][47] ), .A1(out_new[47]), .S(N4740), .Z(n195)
         );
  CMX2X2 U3462 ( .A0(\memory[30][46] ), .A1(out_new[46]), .S(N4740), .Z(n196)
         );
  CMX2X2 U3463 ( .A0(\memory[30][45] ), .A1(out_new[45]), .S(N4740), .Z(n197)
         );
  CMX2X2 U3464 ( .A0(\memory[30][44] ), .A1(out_new[44]), .S(N4740), .Z(n198)
         );
  CMX2X2 U3465 ( .A0(\memory[30][43] ), .A1(out_new[43]), .S(N4740), .Z(n199)
         );
  CMX2X2 U3466 ( .A0(\memory[30][42] ), .A1(out_new[42]), .S(N4740), .Z(n200)
         );
  CMX2X2 U3467 ( .A0(\memory[30][41] ), .A1(out_new[41]), .S(N4740), .Z(n201)
         );
  CMX2X2 U3468 ( .A0(\memory[30][40] ), .A1(out_new[40]), .S(N4740), .Z(n202)
         );
  CMX2X2 U3469 ( .A0(\memory[30][39] ), .A1(out_new[39]), .S(N4740), .Z(n203)
         );
  CMX2X2 U3470 ( .A0(\memory[30][38] ), .A1(out_new[38]), .S(N4740), .Z(n204)
         );
  CMX2X2 U3471 ( .A0(\memory[30][37] ), .A1(out_new[37]), .S(N4740), .Z(n205)
         );
  CMX2X2 U3472 ( .A0(\memory[30][36] ), .A1(out_new[36]), .S(N4740), .Z(n206)
         );
  CMX2X2 U3473 ( .A0(\memory[30][35] ), .A1(out_new[35]), .S(N4740), .Z(n207)
         );
  CMX2X2 U3474 ( .A0(\memory[30][34] ), .A1(out_new[34]), .S(N4740), .Z(n208)
         );
  CMX2X2 U3475 ( .A0(\memory[30][33] ), .A1(out_new[33]), .S(N4740), .Z(n209)
         );
  CMX2X2 U3476 ( .A0(\memory[30][32] ), .A1(out_new[32]), .S(N4740), .Z(n210)
         );
  CMX2X2 U3477 ( .A0(\memory[30][31] ), .A1(out_new[31]), .S(N4740), .Z(n211)
         );
  CMX2X2 U3478 ( .A0(\memory[30][30] ), .A1(out_new[30]), .S(N4740), .Z(n212)
         );
  CMX2X2 U3479 ( .A0(\memory[30][29] ), .A1(out_new[29]), .S(N4740), .Z(n213)
         );
  CMX2X2 U3480 ( .A0(\memory[30][28] ), .A1(out_new[28]), .S(N4740), .Z(n214)
         );
  CMX2X2 U3481 ( .A0(\memory[30][27] ), .A1(out_new[27]), .S(N4740), .Z(n215)
         );
  CMX2X2 U3482 ( .A0(\memory[30][26] ), .A1(out_new[26]), .S(N4740), .Z(n216)
         );
  CMX2X2 U3483 ( .A0(\memory[30][25] ), .A1(out_new[25]), .S(N4740), .Z(n217)
         );
  CMX2X2 U3484 ( .A0(\memory[30][24] ), .A1(out_new[24]), .S(N4740), .Z(n218)
         );
  CMX2X2 U3485 ( .A0(\memory[30][23] ), .A1(out_new[23]), .S(N4740), .Z(n219)
         );
  CMX2X2 U3486 ( .A0(\memory[30][22] ), .A1(out_new[22]), .S(N4740), .Z(n220)
         );
  CMX2X2 U3487 ( .A0(\memory[30][21] ), .A1(out_new[21]), .S(N4740), .Z(n221)
         );
  CMX2X2 U3488 ( .A0(\memory[30][20] ), .A1(out_new[20]), .S(N4740), .Z(n222)
         );
  CMX2X2 U3489 ( .A0(\memory[30][19] ), .A1(out_new[19]), .S(N4740), .Z(n223)
         );
  CMX2X2 U3490 ( .A0(\memory[30][18] ), .A1(out_new[18]), .S(N4740), .Z(n224)
         );
  CMX2X2 U3491 ( .A0(\memory[30][17] ), .A1(out_new[17]), .S(N4740), .Z(n225)
         );
  CMX2X2 U3492 ( .A0(\memory[30][16] ), .A1(out_new[16]), .S(N4740), .Z(n226)
         );
  CMX2X2 U3493 ( .A0(\memory[30][15] ), .A1(out_new[15]), .S(N4740), .Z(n227)
         );
  CMX2X2 U3494 ( .A0(\memory[30][14] ), .A1(out_new[14]), .S(N4740), .Z(n228)
         );
  CMX2X2 U3495 ( .A0(\memory[30][13] ), .A1(out_new[13]), .S(N4740), .Z(n229)
         );
  CMX2X2 U3496 ( .A0(\memory[30][12] ), .A1(out_new[12]), .S(N4740), .Z(n230)
         );
  CMX2X2 U3497 ( .A0(\memory[30][11] ), .A1(out_new[11]), .S(N4740), .Z(n231)
         );
  CMX2X2 U3498 ( .A0(\memory[30][10] ), .A1(out_new[10]), .S(N4740), .Z(n232)
         );
  CMX2X2 U3499 ( .A0(\memory[30][9] ), .A1(out_new[9]), .S(N4740), .Z(n233) );
  CMX2X2 U3500 ( .A0(\memory[30][8] ), .A1(out_new[8]), .S(N4740), .Z(n234) );
  CMX2X2 U3501 ( .A0(\memory[30][7] ), .A1(out_new[7]), .S(N4740), .Z(n235) );
  CMX2X2 U3502 ( .A0(\memory[30][6] ), .A1(out_new[6]), .S(N4740), .Z(n236) );
  CMX2X2 U3503 ( .A0(\memory[30][5] ), .A1(out_new[5]), .S(N4740), .Z(n237) );
  CMX2X2 U3504 ( .A0(\memory[30][4] ), .A1(out_new[4]), .S(N4740), .Z(n238) );
  CMX2X2 U3505 ( .A0(\memory[30][3] ), .A1(out_new[3]), .S(N4740), .Z(n239) );
  CMX2X2 U3506 ( .A0(\memory[30][2] ), .A1(out_new[2]), .S(N4740), .Z(n240) );
  CMX2X2 U3507 ( .A0(\memory[30][1] ), .A1(out_new[1]), .S(N4740), .Z(n241) );
  CMX2X2 U3508 ( .A0(\memory[30][0] ), .A1(out_new[0]), .S(N4740), .Z(n242) );
  CMX2X4 U3509 ( .A0(\memory[29][63] ), .A1(out_new[63]), .S(N4669), .Z(n250)
         );
  CMX2X4 U3510 ( .A0(\memory[29][62] ), .A1(out_new[62]), .S(N4669), .Z(n251)
         );
  CMX2X4 U3511 ( .A0(\memory[29][61] ), .A1(out_new[61]), .S(N4669), .Z(n252)
         );
  CMX2X4 U3512 ( .A0(\memory[29][60] ), .A1(out_new[60]), .S(N4669), .Z(n253)
         );
  CMX2X4 U3513 ( .A0(\memory[29][59] ), .A1(out_new[59]), .S(N4669), .Z(n254)
         );
  CMX2X4 U3514 ( .A0(\memory[29][58] ), .A1(out_new[58]), .S(N4669), .Z(n255)
         );
  CMX2X4 U3515 ( .A0(\memory[29][57] ), .A1(out_new[57]), .S(N4669), .Z(n256)
         );
  CMX2X4 U3516 ( .A0(\memory[29][56] ), .A1(out_new[56]), .S(N4669), .Z(n257)
         );
  CMX2X4 U3517 ( .A0(\memory[29][55] ), .A1(out_new[55]), .S(N4669), .Z(n258)
         );
  CMX2X4 U3518 ( .A0(\memory[29][54] ), .A1(out_new[54]), .S(N4669), .Z(n259)
         );
  CMX2X4 U3519 ( .A0(\memory[29][53] ), .A1(out_new[53]), .S(N4669), .Z(n260)
         );
  CMX2X4 U3520 ( .A0(\memory[29][52] ), .A1(out_new[52]), .S(N4669), .Z(n261)
         );
  CMX2X4 U3521 ( .A0(\memory[29][51] ), .A1(out_new[51]), .S(N4669), .Z(n262)
         );
  CMX2X4 U3522 ( .A0(\memory[29][50] ), .A1(out_new[50]), .S(N4669), .Z(n263)
         );
  CMX2X4 U3523 ( .A0(\memory[29][49] ), .A1(out_new[49]), .S(N4669), .Z(n264)
         );
  CMX2X4 U3524 ( .A0(\memory[29][48] ), .A1(out_new[48]), .S(N4669), .Z(n265)
         );
  CMX2X4 U3525 ( .A0(\memory[29][47] ), .A1(out_new[47]), .S(N4669), .Z(n266)
         );
  CMX2X4 U3526 ( .A0(\memory[29][46] ), .A1(out_new[46]), .S(N4669), .Z(n267)
         );
  CMX2X4 U3527 ( .A0(\memory[29][45] ), .A1(out_new[45]), .S(N4669), .Z(n268)
         );
  CMX2X4 U3528 ( .A0(\memory[29][44] ), .A1(out_new[44]), .S(N4669), .Z(n269)
         );
  CMX2X4 U3529 ( .A0(\memory[29][43] ), .A1(out_new[43]), .S(N4669), .Z(n270)
         );
  CMX2X4 U3530 ( .A0(\memory[29][42] ), .A1(out_new[42]), .S(N4669), .Z(n271)
         );
  CMX2X4 U3531 ( .A0(\memory[29][41] ), .A1(out_new[41]), .S(N4669), .Z(n272)
         );
  CMX2X4 U3532 ( .A0(\memory[29][40] ), .A1(out_new[40]), .S(N4669), .Z(n273)
         );
  CMX2X4 U3533 ( .A0(\memory[29][39] ), .A1(out_new[39]), .S(N4669), .Z(n274)
         );
  CMX2X4 U3534 ( .A0(\memory[29][38] ), .A1(out_new[38]), .S(N4669), .Z(n275)
         );
  CMX2X4 U3535 ( .A0(\memory[29][37] ), .A1(out_new[37]), .S(N4669), .Z(n276)
         );
  CMX2X4 U3536 ( .A0(\memory[29][36] ), .A1(out_new[36]), .S(N4669), .Z(n277)
         );
  CMX2X4 U3537 ( .A0(\memory[29][35] ), .A1(out_new[35]), .S(N4669), .Z(n278)
         );
  CMX2X4 U3538 ( .A0(\memory[29][34] ), .A1(out_new[34]), .S(N4669), .Z(n279)
         );
  CMX2X4 U3539 ( .A0(\memory[29][33] ), .A1(out_new[33]), .S(N4669), .Z(n280)
         );
  CMX2X4 U3540 ( .A0(\memory[29][32] ), .A1(out_new[32]), .S(N4669), .Z(n281)
         );
  CMX2X4 U3541 ( .A0(\memory[29][31] ), .A1(out_new[31]), .S(N4669), .Z(n282)
         );
  CMX2X4 U3542 ( .A0(\memory[29][30] ), .A1(out_new[30]), .S(N4669), .Z(n283)
         );
  CMX2X4 U3543 ( .A0(\memory[29][29] ), .A1(out_new[29]), .S(N4669), .Z(n284)
         );
  CMX2X4 U3544 ( .A0(\memory[29][28] ), .A1(out_new[28]), .S(N4669), .Z(n285)
         );
  CMX2X4 U3545 ( .A0(\memory[29][27] ), .A1(out_new[27]), .S(N4669), .Z(n286)
         );
  CMX2X4 U3546 ( .A0(\memory[29][26] ), .A1(out_new[26]), .S(N4669), .Z(n287)
         );
  CMX2X4 U3547 ( .A0(\memory[29][25] ), .A1(out_new[25]), .S(N4669), .Z(n288)
         );
  CMX2X4 U3548 ( .A0(\memory[29][24] ), .A1(out_new[24]), .S(N4669), .Z(n289)
         );
  CMX2X4 U3549 ( .A0(\memory[29][23] ), .A1(out_new[23]), .S(N4669), .Z(n290)
         );
  CMX2X4 U3550 ( .A0(\memory[29][22] ), .A1(out_new[22]), .S(N4669), .Z(n291)
         );
  CMX2X4 U3551 ( .A0(\memory[29][21] ), .A1(out_new[21]), .S(N4669), .Z(n292)
         );
  CMX2X4 U3552 ( .A0(\memory[29][20] ), .A1(out_new[20]), .S(N4669), .Z(n293)
         );
  CMX2X4 U3553 ( .A0(\memory[29][19] ), .A1(out_new[19]), .S(N4669), .Z(n294)
         );
  CMX2X4 U3554 ( .A0(\memory[29][18] ), .A1(out_new[18]), .S(N4669), .Z(n295)
         );
  CMX2X4 U3555 ( .A0(\memory[29][17] ), .A1(out_new[17]), .S(N4669), .Z(n296)
         );
  CMX2X4 U3556 ( .A0(\memory[29][16] ), .A1(out_new[16]), .S(N4669), .Z(n297)
         );
  CMX2X4 U3557 ( .A0(\memory[29][15] ), .A1(out_new[15]), .S(N4669), .Z(n298)
         );
  CMX2X4 U3558 ( .A0(\memory[29][14] ), .A1(out_new[14]), .S(N4669), .Z(n299)
         );
  CMX2X4 U3559 ( .A0(\memory[29][13] ), .A1(out_new[13]), .S(N4669), .Z(n300)
         );
  CMX2X4 U3560 ( .A0(\memory[29][12] ), .A1(out_new[12]), .S(N4669), .Z(n301)
         );
  CMX2X4 U3561 ( .A0(\memory[29][11] ), .A1(out_new[11]), .S(N4669), .Z(n302)
         );
  CMX2X4 U3562 ( .A0(\memory[29][10] ), .A1(out_new[10]), .S(N4669), .Z(n303)
         );
  CMX2X4 U3563 ( .A0(\memory[29][9] ), .A1(out_new[9]), .S(N4669), .Z(n304) );
  CMX2X4 U3564 ( .A0(\memory[29][8] ), .A1(out_new[8]), .S(N4669), .Z(n305) );
  CMX2X4 U3565 ( .A0(\memory[29][7] ), .A1(out_new[7]), .S(N4669), .Z(n306) );
  CMX2X4 U3566 ( .A0(\memory[29][6] ), .A1(out_new[6]), .S(N4669), .Z(n307) );
  CMX2X4 U3567 ( .A0(\memory[29][5] ), .A1(out_new[5]), .S(N4669), .Z(n308) );
  CMX2X4 U3568 ( .A0(\memory[29][4] ), .A1(out_new[4]), .S(N4669), .Z(n309) );
  CMX2X4 U3569 ( .A0(\memory[29][3] ), .A1(out_new[3]), .S(N4669), .Z(n310) );
  CMX2X4 U3570 ( .A0(\memory[29][2] ), .A1(out_new[2]), .S(N4669), .Z(n311) );
  CMX2X4 U3571 ( .A0(\memory[29][1] ), .A1(out_new[1]), .S(N4669), .Z(n312) );
  CMX2X4 U3572 ( .A0(\memory[29][0] ), .A1(out_new[0]), .S(N4669), .Z(n313) );
  CMX2X2 U3573 ( .A0(\memory[28][63] ), .A1(out_new[63]), .S(N4598), .Z(n321)
         );
  CMX2X2 U3574 ( .A0(\memory[28][62] ), .A1(out_new[62]), .S(N4598), .Z(n322)
         );
  CMX2X2 U3575 ( .A0(\memory[28][61] ), .A1(out_new[61]), .S(N4598), .Z(n323)
         );
  CMX2X2 U3576 ( .A0(\memory[28][60] ), .A1(out_new[60]), .S(N4598), .Z(n324)
         );
  CMX2X2 U3577 ( .A0(\memory[28][59] ), .A1(out_new[59]), .S(N4598), .Z(n325)
         );
  CMX2X2 U3578 ( .A0(\memory[28][58] ), .A1(out_new[58]), .S(N4598), .Z(n326)
         );
  CMX2X2 U3579 ( .A0(\memory[28][57] ), .A1(out_new[57]), .S(N4598), .Z(n327)
         );
  CMX2X2 U3580 ( .A0(\memory[28][56] ), .A1(out_new[56]), .S(N4598), .Z(n328)
         );
  CMX2X2 U3581 ( .A0(\memory[28][55] ), .A1(out_new[55]), .S(N4598), .Z(n329)
         );
  CMX2X2 U3582 ( .A0(\memory[28][54] ), .A1(out_new[54]), .S(N4598), .Z(n330)
         );
  CMX2X2 U3583 ( .A0(\memory[28][53] ), .A1(out_new[53]), .S(N4598), .Z(n331)
         );
  CMX2X2 U3584 ( .A0(\memory[28][52] ), .A1(out_new[52]), .S(N4598), .Z(n332)
         );
  CMX2X2 U3585 ( .A0(\memory[28][51] ), .A1(out_new[51]), .S(N4598), .Z(n333)
         );
  CMX2X2 U3586 ( .A0(\memory[28][50] ), .A1(out_new[50]), .S(N4598), .Z(n334)
         );
  CMX2X2 U3587 ( .A0(\memory[28][49] ), .A1(out_new[49]), .S(N4598), .Z(n335)
         );
  CMX2X2 U3588 ( .A0(\memory[28][48] ), .A1(out_new[48]), .S(N4598), .Z(n336)
         );
  CMX2X2 U3589 ( .A0(\memory[28][47] ), .A1(out_new[47]), .S(N4598), .Z(n337)
         );
  CMX2X2 U3590 ( .A0(\memory[28][46] ), .A1(out_new[46]), .S(N4598), .Z(n338)
         );
  CMX2X2 U3591 ( .A0(\memory[28][45] ), .A1(out_new[45]), .S(N4598), .Z(n339)
         );
  CMX2X2 U3592 ( .A0(\memory[28][44] ), .A1(out_new[44]), .S(N4598), .Z(n340)
         );
  CMX2X2 U3593 ( .A0(\memory[28][43] ), .A1(out_new[43]), .S(N4598), .Z(n341)
         );
  CMX2X2 U3594 ( .A0(\memory[28][42] ), .A1(out_new[42]), .S(N4598), .Z(n342)
         );
  CMX2X2 U3595 ( .A0(\memory[28][41] ), .A1(out_new[41]), .S(N4598), .Z(n343)
         );
  CMX2X2 U3596 ( .A0(\memory[28][40] ), .A1(out_new[40]), .S(N4598), .Z(n344)
         );
  CMX2X2 U3597 ( .A0(\memory[28][39] ), .A1(out_new[39]), .S(N4598), .Z(n345)
         );
  CMX2X2 U3598 ( .A0(\memory[28][38] ), .A1(out_new[38]), .S(N4598), .Z(n346)
         );
  CMX2X2 U3599 ( .A0(\memory[28][37] ), .A1(out_new[37]), .S(N4598), .Z(n347)
         );
  CMX2X2 U3600 ( .A0(\memory[28][36] ), .A1(out_new[36]), .S(N4598), .Z(n348)
         );
  CMX2X2 U3601 ( .A0(\memory[28][35] ), .A1(out_new[35]), .S(N4598), .Z(n349)
         );
  CMX2X2 U3602 ( .A0(\memory[28][34] ), .A1(out_new[34]), .S(N4598), .Z(n350)
         );
  CMX2X2 U3603 ( .A0(\memory[28][33] ), .A1(out_new[33]), .S(N4598), .Z(n351)
         );
  CMX2X2 U3604 ( .A0(\memory[28][32] ), .A1(out_new[32]), .S(N4598), .Z(n352)
         );
  CMX2X2 U3605 ( .A0(\memory[28][31] ), .A1(out_new[31]), .S(N4598), .Z(n353)
         );
  CMX2X2 U3606 ( .A0(\memory[28][30] ), .A1(out_new[30]), .S(N4598), .Z(n354)
         );
  CMX2X2 U3607 ( .A0(\memory[28][29] ), .A1(out_new[29]), .S(N4598), .Z(n355)
         );
  CMX2X2 U3608 ( .A0(\memory[28][28] ), .A1(out_new[28]), .S(N4598), .Z(n356)
         );
  CMX2X2 U3609 ( .A0(\memory[28][27] ), .A1(out_new[27]), .S(N4598), .Z(n357)
         );
  CMX2X2 U3610 ( .A0(\memory[28][26] ), .A1(out_new[26]), .S(N4598), .Z(n358)
         );
  CMX2X2 U3611 ( .A0(\memory[28][25] ), .A1(out_new[25]), .S(N4598), .Z(n359)
         );
  CMX2X2 U3612 ( .A0(\memory[28][24] ), .A1(out_new[24]), .S(N4598), .Z(n360)
         );
  CMX2X2 U3613 ( .A0(\memory[28][23] ), .A1(out_new[23]), .S(N4598), .Z(n361)
         );
  CMX2X2 U3614 ( .A0(\memory[28][22] ), .A1(out_new[22]), .S(N4598), .Z(n362)
         );
  CMX2X2 U3615 ( .A0(\memory[28][21] ), .A1(out_new[21]), .S(N4598), .Z(n363)
         );
  CMX2X2 U3616 ( .A0(\memory[28][20] ), .A1(out_new[20]), .S(N4598), .Z(n364)
         );
  CMX2X2 U3617 ( .A0(\memory[28][19] ), .A1(out_new[19]), .S(N4598), .Z(n365)
         );
  CMX2X2 U3618 ( .A0(\memory[28][18] ), .A1(out_new[18]), .S(N4598), .Z(n366)
         );
  CMX2X2 U3619 ( .A0(\memory[28][17] ), .A1(out_new[17]), .S(N4598), .Z(n367)
         );
  CMX2X2 U3620 ( .A0(\memory[28][16] ), .A1(out_new[16]), .S(N4598), .Z(n368)
         );
  CMX2X2 U3621 ( .A0(\memory[28][15] ), .A1(out_new[15]), .S(N4598), .Z(n369)
         );
  CMX2X2 U3622 ( .A0(\memory[28][14] ), .A1(out_new[14]), .S(N4598), .Z(n370)
         );
  CMX2X2 U3623 ( .A0(\memory[28][13] ), .A1(out_new[13]), .S(N4598), .Z(n371)
         );
  CMX2X2 U3624 ( .A0(\memory[28][12] ), .A1(out_new[12]), .S(N4598), .Z(n372)
         );
  CMX2X2 U3625 ( .A0(\memory[28][11] ), .A1(out_new[11]), .S(N4598), .Z(n373)
         );
  CMX2X2 U3626 ( .A0(\memory[28][10] ), .A1(out_new[10]), .S(N4598), .Z(n374)
         );
  CMX2X2 U3627 ( .A0(\memory[28][9] ), .A1(out_new[9]), .S(N4598), .Z(n375) );
  CMX2X2 U3628 ( .A0(\memory[28][8] ), .A1(out_new[8]), .S(N4598), .Z(n376) );
  CMX2X2 U3629 ( .A0(\memory[28][7] ), .A1(out_new[7]), .S(N4598), .Z(n377) );
  CMX2X2 U3630 ( .A0(\memory[28][6] ), .A1(out_new[6]), .S(N4598), .Z(n378) );
  CMX2X2 U3631 ( .A0(\memory[28][5] ), .A1(out_new[5]), .S(N4598), .Z(n379) );
  CMX2X2 U3632 ( .A0(\memory[28][4] ), .A1(out_new[4]), .S(N4598), .Z(n380) );
  CMX2X2 U3633 ( .A0(\memory[28][3] ), .A1(out_new[3]), .S(N4598), .Z(n381) );
  CMX2X2 U3634 ( .A0(\memory[28][2] ), .A1(out_new[2]), .S(N4598), .Z(n382) );
  CMX2X2 U3635 ( .A0(\memory[28][1] ), .A1(out_new[1]), .S(N4598), .Z(n383) );
  CMX2X2 U3636 ( .A0(\memory[28][0] ), .A1(out_new[0]), .S(N4598), .Z(n384) );
  CMX2X2 U3637 ( .A0(\memory[26][63] ), .A1(out_new[63]), .S(N4456), .Z(n463)
         );
  CMX2X2 U3638 ( .A0(\memory[26][62] ), .A1(out_new[62]), .S(N4456), .Z(n464)
         );
  CMX2X2 U3639 ( .A0(\memory[26][61] ), .A1(out_new[61]), .S(N4456), .Z(n465)
         );
  CMX2X2 U3640 ( .A0(\memory[26][60] ), .A1(out_new[60]), .S(N4456), .Z(n466)
         );
  CMX2X2 U3641 ( .A0(\memory[26][59] ), .A1(out_new[59]), .S(N4456), .Z(n467)
         );
  CMX2X2 U3642 ( .A0(\memory[26][58] ), .A1(out_new[58]), .S(N4456), .Z(n468)
         );
  CMX2X2 U3643 ( .A0(\memory[26][57] ), .A1(out_new[57]), .S(N4456), .Z(n469)
         );
  CMX2X2 U3644 ( .A0(\memory[26][56] ), .A1(out_new[56]), .S(N4456), .Z(n470)
         );
  CMX2X2 U3645 ( .A0(\memory[26][55] ), .A1(out_new[55]), .S(N4456), .Z(n471)
         );
  CMX2X2 U3646 ( .A0(\memory[26][54] ), .A1(out_new[54]), .S(N4456), .Z(n472)
         );
  CMX2X2 U3647 ( .A0(\memory[26][53] ), .A1(out_new[53]), .S(N4456), .Z(n473)
         );
  CMX2X2 U3648 ( .A0(\memory[26][52] ), .A1(out_new[52]), .S(N4456), .Z(n474)
         );
  CMX2X2 U3649 ( .A0(\memory[26][51] ), .A1(out_new[51]), .S(N4456), .Z(n475)
         );
  CMX2X2 U3650 ( .A0(\memory[26][50] ), .A1(out_new[50]), .S(N4456), .Z(n476)
         );
  CMX2X2 U3651 ( .A0(\memory[26][49] ), .A1(out_new[49]), .S(N4456), .Z(n477)
         );
  CMX2X2 U3652 ( .A0(\memory[26][48] ), .A1(out_new[48]), .S(N4456), .Z(n478)
         );
  CMX2X2 U3653 ( .A0(\memory[26][47] ), .A1(out_new[47]), .S(N4456), .Z(n479)
         );
  CMX2X2 U3654 ( .A0(\memory[26][46] ), .A1(out_new[46]), .S(N4456), .Z(n480)
         );
  CMX2X2 U3655 ( .A0(\memory[26][45] ), .A1(out_new[45]), .S(N4456), .Z(n481)
         );
  CMX2X2 U3656 ( .A0(\memory[26][44] ), .A1(out_new[44]), .S(N4456), .Z(n482)
         );
  CMX2X2 U3657 ( .A0(\memory[26][43] ), .A1(out_new[43]), .S(N4456), .Z(n483)
         );
  CMX2X2 U3658 ( .A0(\memory[26][42] ), .A1(out_new[42]), .S(N4456), .Z(n484)
         );
  CMX2X2 U3659 ( .A0(\memory[26][41] ), .A1(out_new[41]), .S(N4456), .Z(n485)
         );
  CMX2X2 U3660 ( .A0(\memory[26][40] ), .A1(out_new[40]), .S(N4456), .Z(n486)
         );
  CMX2X2 U3661 ( .A0(\memory[26][39] ), .A1(out_new[39]), .S(N4456), .Z(n487)
         );
  CMX2X2 U3662 ( .A0(\memory[26][38] ), .A1(out_new[38]), .S(N4456), .Z(n488)
         );
  CMX2X2 U3663 ( .A0(\memory[26][37] ), .A1(out_new[37]), .S(N4456), .Z(n489)
         );
  CMX2X2 U3664 ( .A0(\memory[26][36] ), .A1(out_new[36]), .S(N4456), .Z(n490)
         );
  CMX2X2 U3665 ( .A0(\memory[26][35] ), .A1(out_new[35]), .S(N4456), .Z(n491)
         );
  CMX2X2 U3666 ( .A0(\memory[26][34] ), .A1(out_new[34]), .S(N4456), .Z(n492)
         );
  CMX2X2 U3667 ( .A0(\memory[26][33] ), .A1(out_new[33]), .S(N4456), .Z(n493)
         );
  CMX2X2 U3668 ( .A0(\memory[26][32] ), .A1(out_new[32]), .S(N4456), .Z(n494)
         );
  CMX2X2 U3669 ( .A0(\memory[26][31] ), .A1(out_new[31]), .S(N4456), .Z(n495)
         );
  CMX2X2 U3670 ( .A0(\memory[26][30] ), .A1(out_new[30]), .S(N4456), .Z(n496)
         );
  CMX2X2 U3671 ( .A0(\memory[26][29] ), .A1(out_new[29]), .S(N4456), .Z(n497)
         );
  CMX2X2 U3672 ( .A0(\memory[26][28] ), .A1(out_new[28]), .S(N4456), .Z(n498)
         );
  CMX2X2 U3673 ( .A0(\memory[26][27] ), .A1(out_new[27]), .S(N4456), .Z(n499)
         );
  CMX2X2 U3674 ( .A0(\memory[26][26] ), .A1(out_new[26]), .S(N4456), .Z(n500)
         );
  CMX2X2 U3675 ( .A0(\memory[26][25] ), .A1(out_new[25]), .S(N4456), .Z(n501)
         );
  CMX2X2 U3676 ( .A0(\memory[26][24] ), .A1(out_new[24]), .S(N4456), .Z(n502)
         );
  CMX2X2 U3677 ( .A0(\memory[26][23] ), .A1(out_new[23]), .S(N4456), .Z(n503)
         );
  CMX2X2 U3678 ( .A0(\memory[26][22] ), .A1(out_new[22]), .S(N4456), .Z(n504)
         );
  CMX2X2 U3679 ( .A0(\memory[26][21] ), .A1(out_new[21]), .S(N4456), .Z(n505)
         );
  CMX2X2 U3680 ( .A0(\memory[26][20] ), .A1(out_new[20]), .S(N4456), .Z(n506)
         );
  CMX2X2 U3681 ( .A0(\memory[26][19] ), .A1(out_new[19]), .S(N4456), .Z(n507)
         );
  CMX2X2 U3682 ( .A0(\memory[26][18] ), .A1(out_new[18]), .S(N4456), .Z(n508)
         );
  CMX2X2 U3683 ( .A0(\memory[26][17] ), .A1(out_new[17]), .S(N4456), .Z(n509)
         );
  CMX2X2 U3684 ( .A0(\memory[26][16] ), .A1(out_new[16]), .S(N4456), .Z(n510)
         );
  CMX2X2 U3685 ( .A0(\memory[26][15] ), .A1(out_new[15]), .S(N4456), .Z(n511)
         );
  CMX2X2 U3686 ( .A0(\memory[26][14] ), .A1(out_new[14]), .S(N4456), .Z(n512)
         );
  CMX2X2 U3687 ( .A0(\memory[26][13] ), .A1(out_new[13]), .S(N4456), .Z(n513)
         );
  CMX2X2 U3688 ( .A0(\memory[26][12] ), .A1(out_new[12]), .S(N4456), .Z(n514)
         );
  CMX2X2 U3689 ( .A0(\memory[26][11] ), .A1(out_new[11]), .S(N4456), .Z(n515)
         );
  CMX2X2 U3690 ( .A0(\memory[26][10] ), .A1(out_new[10]), .S(N4456), .Z(n516)
         );
  CMX2X2 U3691 ( .A0(\memory[26][9] ), .A1(out_new[9]), .S(N4456), .Z(n517) );
  CMX2X2 U3692 ( .A0(\memory[26][8] ), .A1(out_new[8]), .S(N4456), .Z(n518) );
  CMX2X2 U3693 ( .A0(\memory[26][7] ), .A1(out_new[7]), .S(N4456), .Z(n519) );
  CMX2X2 U3694 ( .A0(\memory[26][6] ), .A1(out_new[6]), .S(N4456), .Z(n520) );
  CMX2X2 U3695 ( .A0(\memory[26][5] ), .A1(out_new[5]), .S(N4456), .Z(n521) );
  CMX2X2 U3696 ( .A0(\memory[26][4] ), .A1(out_new[4]), .S(N4456), .Z(n522) );
  CMX2X2 U3697 ( .A0(\memory[26][3] ), .A1(out_new[3]), .S(N4456), .Z(n523) );
  CMX2X2 U3698 ( .A0(\memory[26][2] ), .A1(out_new[2]), .S(N4456), .Z(n524) );
  CMX2X2 U3699 ( .A0(\memory[26][1] ), .A1(out_new[1]), .S(N4456), .Z(n525) );
  CMX2X2 U3700 ( .A0(\memory[26][0] ), .A1(out_new[0]), .S(N4456), .Z(n526) );
  CMX2X2 U3701 ( .A0(\memory[25][63] ), .A1(out_new[63]), .S(N4385), .Z(n534)
         );
  CMX2X2 U3702 ( .A0(\memory[25][62] ), .A1(out_new[62]), .S(N4385), .Z(n535)
         );
  CMX2X2 U3703 ( .A0(\memory[25][61] ), .A1(out_new[61]), .S(N4385), .Z(n536)
         );
  CMX2X2 U3704 ( .A0(\memory[25][60] ), .A1(out_new[60]), .S(N4385), .Z(n537)
         );
  CMX2X2 U3705 ( .A0(\memory[25][59] ), .A1(out_new[59]), .S(N4385), .Z(n538)
         );
  CMX2X2 U3706 ( .A0(\memory[25][58] ), .A1(out_new[58]), .S(N4385), .Z(n539)
         );
  CMX2X2 U3707 ( .A0(\memory[25][57] ), .A1(out_new[57]), .S(N4385), .Z(n540)
         );
  CMX2X2 U3708 ( .A0(\memory[25][56] ), .A1(out_new[56]), .S(N4385), .Z(n541)
         );
  CMX2X2 U3709 ( .A0(\memory[25][55] ), .A1(out_new[55]), .S(N4385), .Z(n542)
         );
  CMX2X2 U3710 ( .A0(\memory[25][54] ), .A1(out_new[54]), .S(N4385), .Z(n543)
         );
  CMX2X2 U3711 ( .A0(\memory[25][53] ), .A1(out_new[53]), .S(N4385), .Z(n544)
         );
  CMX2X2 U3712 ( .A0(\memory[25][52] ), .A1(out_new[52]), .S(N4385), .Z(n545)
         );
  CMX2X2 U3713 ( .A0(\memory[25][51] ), .A1(out_new[51]), .S(N4385), .Z(n546)
         );
  CMX2X2 U3714 ( .A0(\memory[25][50] ), .A1(out_new[50]), .S(N4385), .Z(n547)
         );
  CMX2X2 U3715 ( .A0(\memory[25][49] ), .A1(out_new[49]), .S(N4385), .Z(n548)
         );
  CMX2X2 U3716 ( .A0(\memory[25][48] ), .A1(out_new[48]), .S(N4385), .Z(n549)
         );
  CMX2X2 U3717 ( .A0(\memory[25][47] ), .A1(out_new[47]), .S(N4385), .Z(n550)
         );
  CMX2X2 U3718 ( .A0(\memory[25][46] ), .A1(out_new[46]), .S(N4385), .Z(n551)
         );
  CMX2X2 U3719 ( .A0(\memory[25][45] ), .A1(out_new[45]), .S(N4385), .Z(n552)
         );
  CMX2X2 U3720 ( .A0(\memory[25][44] ), .A1(out_new[44]), .S(N4385), .Z(n553)
         );
  CMX2X2 U3721 ( .A0(\memory[25][43] ), .A1(out_new[43]), .S(N4385), .Z(n554)
         );
  CMX2X2 U3722 ( .A0(\memory[25][42] ), .A1(out_new[42]), .S(N4385), .Z(n555)
         );
  CMX2X2 U3723 ( .A0(\memory[25][41] ), .A1(out_new[41]), .S(N4385), .Z(n556)
         );
  CMX2X2 U3724 ( .A0(\memory[25][40] ), .A1(out_new[40]), .S(N4385), .Z(n557)
         );
  CMX2X2 U3725 ( .A0(\memory[25][39] ), .A1(out_new[39]), .S(N4385), .Z(n558)
         );
  CMX2X2 U3726 ( .A0(\memory[25][38] ), .A1(out_new[38]), .S(N4385), .Z(n559)
         );
  CMX2X2 U3727 ( .A0(\memory[25][37] ), .A1(out_new[37]), .S(N4385), .Z(n560)
         );
  CMX2X2 U3728 ( .A0(\memory[25][36] ), .A1(out_new[36]), .S(N4385), .Z(n561)
         );
  CMX2X2 U3729 ( .A0(\memory[25][35] ), .A1(out_new[35]), .S(N4385), .Z(n562)
         );
  CMX2X2 U3730 ( .A0(\memory[25][34] ), .A1(out_new[34]), .S(N4385), .Z(n563)
         );
  CMX2X2 U3731 ( .A0(\memory[25][33] ), .A1(out_new[33]), .S(N4385), .Z(n564)
         );
  CMX2X2 U3732 ( .A0(\memory[25][32] ), .A1(out_new[32]), .S(N4385), .Z(n565)
         );
  CMX2X2 U3733 ( .A0(\memory[25][31] ), .A1(out_new[31]), .S(N4385), .Z(n566)
         );
  CMX2X2 U3734 ( .A0(\memory[25][30] ), .A1(out_new[30]), .S(N4385), .Z(n567)
         );
  CMX2X2 U3735 ( .A0(\memory[25][29] ), .A1(out_new[29]), .S(N4385), .Z(n568)
         );
  CMX2X2 U3736 ( .A0(\memory[25][28] ), .A1(out_new[28]), .S(N4385), .Z(n569)
         );
  CMX2X2 U3737 ( .A0(\memory[25][27] ), .A1(out_new[27]), .S(N4385), .Z(n570)
         );
  CMX2X2 U3738 ( .A0(\memory[25][26] ), .A1(out_new[26]), .S(N4385), .Z(n571)
         );
  CMX2X2 U3739 ( .A0(\memory[25][25] ), .A1(out_new[25]), .S(N4385), .Z(n572)
         );
  CMX2X2 U3740 ( .A0(\memory[25][24] ), .A1(out_new[24]), .S(N4385), .Z(n573)
         );
  CMX2X2 U3741 ( .A0(\memory[25][23] ), .A1(out_new[23]), .S(N4385), .Z(n574)
         );
  CMX2X2 U3742 ( .A0(\memory[25][22] ), .A1(out_new[22]), .S(N4385), .Z(n575)
         );
  CMX2X2 U3743 ( .A0(\memory[25][21] ), .A1(out_new[21]), .S(N4385), .Z(n576)
         );
  CMX2X2 U3744 ( .A0(\memory[25][20] ), .A1(out_new[20]), .S(N4385), .Z(n577)
         );
  CMX2X2 U3745 ( .A0(\memory[25][19] ), .A1(out_new[19]), .S(N4385), .Z(n578)
         );
  CMX2X2 U3746 ( .A0(\memory[25][18] ), .A1(out_new[18]), .S(N4385), .Z(n579)
         );
  CMX2X2 U3747 ( .A0(\memory[25][17] ), .A1(out_new[17]), .S(N4385), .Z(n580)
         );
  CMX2X2 U3748 ( .A0(\memory[25][16] ), .A1(out_new[16]), .S(N4385), .Z(n581)
         );
  CMX2X2 U3749 ( .A0(\memory[25][15] ), .A1(out_new[15]), .S(N4385), .Z(n582)
         );
  CMX2X2 U3750 ( .A0(\memory[25][14] ), .A1(out_new[14]), .S(N4385), .Z(n583)
         );
  CMX2X2 U3751 ( .A0(\memory[25][13] ), .A1(out_new[13]), .S(N4385), .Z(n584)
         );
  CMX2X2 U3752 ( .A0(\memory[25][12] ), .A1(out_new[12]), .S(N4385), .Z(n585)
         );
  CMX2X2 U3753 ( .A0(\memory[25][11] ), .A1(out_new[11]), .S(N4385), .Z(n586)
         );
  CMX2X2 U3754 ( .A0(\memory[25][10] ), .A1(out_new[10]), .S(N4385), .Z(n587)
         );
  CMX2X2 U3755 ( .A0(\memory[25][9] ), .A1(out_new[9]), .S(N4385), .Z(n588) );
  CMX2X2 U3756 ( .A0(\memory[25][8] ), .A1(out_new[8]), .S(N4385), .Z(n589) );
  CMX2X2 U3757 ( .A0(\memory[25][7] ), .A1(out_new[7]), .S(N4385), .Z(n590) );
  CMX2X2 U3758 ( .A0(\memory[25][6] ), .A1(out_new[6]), .S(N4385), .Z(n591) );
  CMX2X2 U3759 ( .A0(\memory[25][5] ), .A1(out_new[5]), .S(N4385), .Z(n592) );
  CMX2X2 U3760 ( .A0(\memory[25][4] ), .A1(out_new[4]), .S(N4385), .Z(n593) );
  CMX2X2 U3761 ( .A0(\memory[25][3] ), .A1(out_new[3]), .S(N4385), .Z(n594) );
  CMX2X2 U3762 ( .A0(\memory[25][2] ), .A1(out_new[2]), .S(N4385), .Z(n595) );
  CMX2X2 U3763 ( .A0(\memory[25][1] ), .A1(out_new[1]), .S(N4385), .Z(n596) );
  CMX2X2 U3764 ( .A0(\memory[25][0] ), .A1(out_new[0]), .S(N4385), .Z(n597) );
  CMX2X2 U3765 ( .A0(\memory[24][63] ), .A1(out_new[63]), .S(N4314), .Z(n605)
         );
  CMX2X2 U3766 ( .A0(\memory[24][62] ), .A1(out_new[62]), .S(N4314), .Z(n606)
         );
  CMX2X2 U3767 ( .A0(\memory[24][61] ), .A1(out_new[61]), .S(N4314), .Z(n607)
         );
  CMX2X2 U3768 ( .A0(\memory[24][60] ), .A1(out_new[60]), .S(N4314), .Z(n608)
         );
  CMX2X2 U3769 ( .A0(\memory[24][59] ), .A1(out_new[59]), .S(N4314), .Z(n609)
         );
  CMX2X2 U3770 ( .A0(\memory[24][58] ), .A1(out_new[58]), .S(N4314), .Z(n610)
         );
  CMX2X2 U3771 ( .A0(\memory[24][57] ), .A1(out_new[57]), .S(N4314), .Z(n611)
         );
  CMX2X2 U3772 ( .A0(\memory[24][56] ), .A1(out_new[56]), .S(N4314), .Z(n612)
         );
  CMX2X2 U3773 ( .A0(\memory[24][55] ), .A1(out_new[55]), .S(N4314), .Z(n613)
         );
  CMX2X2 U3774 ( .A0(\memory[24][54] ), .A1(out_new[54]), .S(N4314), .Z(n614)
         );
  CMX2X2 U3775 ( .A0(\memory[24][53] ), .A1(out_new[53]), .S(N4314), .Z(n615)
         );
  CMX2X2 U3776 ( .A0(\memory[24][52] ), .A1(out_new[52]), .S(N4314), .Z(n616)
         );
  CMX2X2 U3777 ( .A0(\memory[24][51] ), .A1(out_new[51]), .S(N4314), .Z(n617)
         );
  CMX2X2 U3778 ( .A0(\memory[24][50] ), .A1(out_new[50]), .S(N4314), .Z(n618)
         );
  CMX2X2 U3779 ( .A0(\memory[24][49] ), .A1(out_new[49]), .S(N4314), .Z(n619)
         );
  CMX2X2 U3780 ( .A0(\memory[24][48] ), .A1(out_new[48]), .S(N4314), .Z(n620)
         );
  CMX2X2 U3781 ( .A0(\memory[24][47] ), .A1(out_new[47]), .S(N4314), .Z(n621)
         );
  CMX2X2 U3782 ( .A0(\memory[24][46] ), .A1(out_new[46]), .S(N4314), .Z(n622)
         );
  CMX2X2 U3783 ( .A0(\memory[24][45] ), .A1(out_new[45]), .S(N4314), .Z(n623)
         );
  CMX2X2 U3784 ( .A0(\memory[24][44] ), .A1(out_new[44]), .S(N4314), .Z(n624)
         );
  CMX2X2 U3785 ( .A0(\memory[24][43] ), .A1(out_new[43]), .S(N4314), .Z(n625)
         );
  CMX2X2 U3786 ( .A0(\memory[24][42] ), .A1(out_new[42]), .S(N4314), .Z(n626)
         );
  CMX2X2 U3787 ( .A0(\memory[24][41] ), .A1(out_new[41]), .S(N4314), .Z(n627)
         );
  CMX2X2 U3788 ( .A0(\memory[24][40] ), .A1(out_new[40]), .S(N4314), .Z(n628)
         );
  CMX2X2 U3789 ( .A0(\memory[24][39] ), .A1(out_new[39]), .S(N4314), .Z(n629)
         );
  CMX2X2 U3790 ( .A0(\memory[24][38] ), .A1(out_new[38]), .S(N4314), .Z(n630)
         );
  CMX2X2 U3791 ( .A0(\memory[24][37] ), .A1(out_new[37]), .S(N4314), .Z(n631)
         );
  CMX2X2 U3792 ( .A0(\memory[24][36] ), .A1(out_new[36]), .S(N4314), .Z(n632)
         );
  CMX2X2 U3793 ( .A0(\memory[24][35] ), .A1(out_new[35]), .S(N4314), .Z(n633)
         );
  CMX2X2 U3794 ( .A0(\memory[24][34] ), .A1(out_new[34]), .S(N4314), .Z(n634)
         );
  CMX2X2 U3795 ( .A0(\memory[24][33] ), .A1(out_new[33]), .S(N4314), .Z(n635)
         );
  CMX2X2 U3796 ( .A0(\memory[24][32] ), .A1(out_new[32]), .S(N4314), .Z(n636)
         );
  CMX2X2 U3797 ( .A0(\memory[24][31] ), .A1(out_new[31]), .S(N4314), .Z(n637)
         );
  CMX2X2 U3798 ( .A0(\memory[24][30] ), .A1(out_new[30]), .S(N4314), .Z(n638)
         );
  CMX2X2 U3799 ( .A0(\memory[24][29] ), .A1(out_new[29]), .S(N4314), .Z(n639)
         );
  CMX2X2 U3800 ( .A0(\memory[24][28] ), .A1(out_new[28]), .S(N4314), .Z(n640)
         );
  CMX2X2 U3801 ( .A0(\memory[24][27] ), .A1(out_new[27]), .S(N4314), .Z(n641)
         );
  CMX2X2 U3802 ( .A0(\memory[24][26] ), .A1(out_new[26]), .S(N4314), .Z(n642)
         );
  CMX2X2 U3803 ( .A0(\memory[24][25] ), .A1(out_new[25]), .S(N4314), .Z(n643)
         );
  CMX2X2 U3804 ( .A0(\memory[24][24] ), .A1(out_new[24]), .S(N4314), .Z(n644)
         );
  CMX2X2 U3805 ( .A0(\memory[24][23] ), .A1(out_new[23]), .S(N4314), .Z(n645)
         );
  CMX2X2 U3806 ( .A0(\memory[24][22] ), .A1(out_new[22]), .S(N4314), .Z(n646)
         );
  CMX2X2 U3807 ( .A0(\memory[24][21] ), .A1(out_new[21]), .S(N4314), .Z(n647)
         );
  CMX2X2 U3808 ( .A0(\memory[24][20] ), .A1(out_new[20]), .S(N4314), .Z(n648)
         );
  CMX2X2 U3809 ( .A0(\memory[24][19] ), .A1(out_new[19]), .S(N4314), .Z(n649)
         );
  CMX2X2 U3810 ( .A0(\memory[24][18] ), .A1(out_new[18]), .S(N4314), .Z(n650)
         );
  CMX2X2 U3811 ( .A0(\memory[24][17] ), .A1(out_new[17]), .S(N4314), .Z(n651)
         );
  CMX2X2 U3812 ( .A0(\memory[24][16] ), .A1(out_new[16]), .S(N4314), .Z(n652)
         );
  CMX2X2 U3813 ( .A0(\memory[24][15] ), .A1(out_new[15]), .S(N4314), .Z(n653)
         );
  CMX2X2 U3814 ( .A0(\memory[24][14] ), .A1(out_new[14]), .S(N4314), .Z(n654)
         );
  CMX2X2 U3815 ( .A0(\memory[24][13] ), .A1(out_new[13]), .S(N4314), .Z(n655)
         );
  CMX2X2 U3816 ( .A0(\memory[24][12] ), .A1(out_new[12]), .S(N4314), .Z(n656)
         );
  CMX2X2 U3817 ( .A0(\memory[24][11] ), .A1(out_new[11]), .S(N4314), .Z(n657)
         );
  CMX2X2 U3818 ( .A0(\memory[24][10] ), .A1(out_new[10]), .S(N4314), .Z(n658)
         );
  CMX2X2 U3819 ( .A0(\memory[24][9] ), .A1(out_new[9]), .S(N4314), .Z(n659) );
  CMX2X2 U3820 ( .A0(\memory[24][8] ), .A1(out_new[8]), .S(N4314), .Z(n660) );
  CMX2X2 U3821 ( .A0(\memory[24][7] ), .A1(out_new[7]), .S(N4314), .Z(n661) );
  CMX2X2 U3822 ( .A0(\memory[24][6] ), .A1(out_new[6]), .S(N4314), .Z(n662) );
  CMX2X2 U3823 ( .A0(\memory[24][5] ), .A1(out_new[5]), .S(N4314), .Z(n663) );
  CMX2X2 U3824 ( .A0(\memory[24][4] ), .A1(out_new[4]), .S(N4314), .Z(n664) );
  CMX2X2 U3825 ( .A0(\memory[24][3] ), .A1(out_new[3]), .S(N4314), .Z(n665) );
  CMX2X2 U3826 ( .A0(\memory[24][2] ), .A1(out_new[2]), .S(N4314), .Z(n666) );
  CMX2X2 U3827 ( .A0(\memory[24][1] ), .A1(out_new[1]), .S(N4314), .Z(n667) );
  CMX2X2 U3828 ( .A0(\memory[24][0] ), .A1(out_new[0]), .S(N4314), .Z(n668) );
  CMX2X2 U3829 ( .A0(\memory[22][63] ), .A1(out_new[63]), .S(N4172), .Z(n747)
         );
  CMX2X2 U3830 ( .A0(\memory[22][62] ), .A1(out_new[62]), .S(N4172), .Z(n748)
         );
  CMX2X2 U3831 ( .A0(\memory[22][61] ), .A1(out_new[61]), .S(N4172), .Z(n749)
         );
  CMX2X2 U3832 ( .A0(\memory[22][60] ), .A1(out_new[60]), .S(N4172), .Z(n750)
         );
  CMX2X2 U3833 ( .A0(\memory[22][59] ), .A1(out_new[59]), .S(N4172), .Z(n751)
         );
  CMX2X2 U3834 ( .A0(\memory[22][58] ), .A1(out_new[58]), .S(N4172), .Z(n752)
         );
  CMX2X2 U3835 ( .A0(\memory[22][57] ), .A1(out_new[57]), .S(N4172), .Z(n753)
         );
  CMX2X2 U3836 ( .A0(\memory[22][56] ), .A1(out_new[56]), .S(N4172), .Z(n754)
         );
  CMX2X2 U3837 ( .A0(\memory[22][55] ), .A1(out_new[55]), .S(N4172), .Z(n755)
         );
  CMX2X2 U3838 ( .A0(\memory[22][54] ), .A1(out_new[54]), .S(N4172), .Z(n756)
         );
  CMX2X2 U3839 ( .A0(\memory[22][53] ), .A1(out_new[53]), .S(N4172), .Z(n757)
         );
  CMX2X2 U3840 ( .A0(\memory[22][52] ), .A1(out_new[52]), .S(N4172), .Z(n758)
         );
  CMX2X2 U3841 ( .A0(\memory[22][51] ), .A1(out_new[51]), .S(N4172), .Z(n759)
         );
  CMX2X2 U3842 ( .A0(\memory[22][50] ), .A1(out_new[50]), .S(N4172), .Z(n760)
         );
  CMX2X2 U3843 ( .A0(\memory[22][49] ), .A1(out_new[49]), .S(N4172), .Z(n761)
         );
  CMX2X2 U3844 ( .A0(\memory[22][48] ), .A1(out_new[48]), .S(N4172), .Z(n762)
         );
  CMX2X2 U3845 ( .A0(\memory[22][47] ), .A1(out_new[47]), .S(N4172), .Z(n763)
         );
  CMX2X2 U3846 ( .A0(\memory[22][46] ), .A1(out_new[46]), .S(N4172), .Z(n764)
         );
  CMX2X2 U3847 ( .A0(\memory[22][45] ), .A1(out_new[45]), .S(N4172), .Z(n765)
         );
  CMX2X2 U3848 ( .A0(\memory[22][44] ), .A1(out_new[44]), .S(N4172), .Z(n766)
         );
  CMX2X2 U3849 ( .A0(\memory[22][43] ), .A1(out_new[43]), .S(N4172), .Z(n767)
         );
  CMX2X2 U3850 ( .A0(\memory[22][42] ), .A1(out_new[42]), .S(N4172), .Z(n768)
         );
  CMX2X2 U3851 ( .A0(\memory[22][41] ), .A1(out_new[41]), .S(N4172), .Z(n769)
         );
  CMX2X2 U3852 ( .A0(\memory[22][40] ), .A1(out_new[40]), .S(N4172), .Z(n770)
         );
  CMX2X2 U3853 ( .A0(\memory[22][39] ), .A1(out_new[39]), .S(N4172), .Z(n771)
         );
  CMX2X2 U3854 ( .A0(\memory[22][38] ), .A1(out_new[38]), .S(N4172), .Z(n772)
         );
  CMX2X2 U3855 ( .A0(\memory[22][37] ), .A1(out_new[37]), .S(N4172), .Z(n773)
         );
  CMX2X2 U3856 ( .A0(\memory[22][36] ), .A1(out_new[36]), .S(N4172), .Z(n774)
         );
  CMX2X2 U3857 ( .A0(\memory[22][35] ), .A1(out_new[35]), .S(N4172), .Z(n775)
         );
  CMX2X2 U3858 ( .A0(\memory[22][34] ), .A1(out_new[34]), .S(N4172), .Z(n776)
         );
  CMX2X2 U3859 ( .A0(\memory[22][33] ), .A1(out_new[33]), .S(N4172), .Z(n777)
         );
  CMX2X2 U3860 ( .A0(\memory[22][32] ), .A1(out_new[32]), .S(N4172), .Z(n778)
         );
  CMX2X2 U3861 ( .A0(\memory[22][31] ), .A1(out_new[31]), .S(N4172), .Z(n779)
         );
  CMX2X2 U3862 ( .A0(\memory[22][30] ), .A1(out_new[30]), .S(N4172), .Z(n780)
         );
  CMX2X2 U3863 ( .A0(\memory[22][29] ), .A1(out_new[29]), .S(N4172), .Z(n781)
         );
  CMX2X2 U3864 ( .A0(\memory[22][28] ), .A1(out_new[28]), .S(N4172), .Z(n782)
         );
  CMX2X2 U3865 ( .A0(\memory[22][27] ), .A1(out_new[27]), .S(N4172), .Z(n783)
         );
  CMX2X2 U3866 ( .A0(\memory[22][26] ), .A1(out_new[26]), .S(N4172), .Z(n784)
         );
  CMX2X2 U3867 ( .A0(\memory[22][25] ), .A1(out_new[25]), .S(N4172), .Z(n785)
         );
  CMX2X2 U3868 ( .A0(\memory[22][24] ), .A1(out_new[24]), .S(N4172), .Z(n786)
         );
  CMX2X2 U3869 ( .A0(\memory[22][23] ), .A1(out_new[23]), .S(N4172), .Z(n787)
         );
  CMX2X2 U3870 ( .A0(\memory[22][22] ), .A1(out_new[22]), .S(N4172), .Z(n788)
         );
  CMX2X2 U3871 ( .A0(\memory[22][21] ), .A1(out_new[21]), .S(N4172), .Z(n789)
         );
  CMX2X2 U3872 ( .A0(\memory[22][20] ), .A1(out_new[20]), .S(N4172), .Z(n790)
         );
  CMX2X2 U3873 ( .A0(\memory[22][19] ), .A1(out_new[19]), .S(N4172), .Z(n791)
         );
  CMX2X2 U3874 ( .A0(\memory[22][18] ), .A1(out_new[18]), .S(N4172), .Z(n792)
         );
  CMX2X2 U3875 ( .A0(\memory[22][17] ), .A1(out_new[17]), .S(N4172), .Z(n793)
         );
  CMX2X2 U3876 ( .A0(\memory[22][16] ), .A1(out_new[16]), .S(N4172), .Z(n794)
         );
  CMX2X2 U3877 ( .A0(\memory[22][15] ), .A1(out_new[15]), .S(N4172), .Z(n795)
         );
  CMX2X2 U3878 ( .A0(\memory[22][14] ), .A1(out_new[14]), .S(N4172), .Z(n796)
         );
  CMX2X2 U3879 ( .A0(\memory[22][13] ), .A1(out_new[13]), .S(N4172), .Z(n797)
         );
  CMX2X2 U3880 ( .A0(\memory[22][12] ), .A1(out_new[12]), .S(N4172), .Z(n798)
         );
  CMX2X2 U3881 ( .A0(\memory[22][11] ), .A1(out_new[11]), .S(N4172), .Z(n799)
         );
  CMX2X2 U3882 ( .A0(\memory[22][10] ), .A1(out_new[10]), .S(N4172), .Z(n800)
         );
  CMX2X2 U3883 ( .A0(\memory[22][9] ), .A1(out_new[9]), .S(N4172), .Z(n801) );
  CMX2X2 U3884 ( .A0(\memory[22][8] ), .A1(out_new[8]), .S(N4172), .Z(n802) );
  CMX2X2 U3885 ( .A0(\memory[22][7] ), .A1(out_new[7]), .S(N4172), .Z(n803) );
  CMX2X2 U3886 ( .A0(\memory[22][6] ), .A1(out_new[6]), .S(N4172), .Z(n804) );
  CMX2X2 U3887 ( .A0(\memory[22][5] ), .A1(out_new[5]), .S(N4172), .Z(n805) );
  CMX2X2 U3888 ( .A0(\memory[22][4] ), .A1(out_new[4]), .S(N4172), .Z(n806) );
  CMX2X2 U3889 ( .A0(\memory[22][3] ), .A1(out_new[3]), .S(N4172), .Z(n807) );
  CMX2X2 U3890 ( .A0(\memory[22][2] ), .A1(out_new[2]), .S(N4172), .Z(n808) );
  CMX2X2 U3891 ( .A0(\memory[22][1] ), .A1(out_new[1]), .S(N4172), .Z(n809) );
  CMX2X2 U3892 ( .A0(\memory[22][0] ), .A1(out_new[0]), .S(N4172), .Z(n810) );
  CMX2X4 U3893 ( .A0(\memory[21][63] ), .A1(out_new[63]), .S(N4101), .Z(n818)
         );
  CMX2X4 U3894 ( .A0(\memory[21][62] ), .A1(out_new[62]), .S(N4101), .Z(n819)
         );
  CMX2X4 U3895 ( .A0(\memory[21][61] ), .A1(out_new[61]), .S(N4101), .Z(n820)
         );
  CMX2X4 U3896 ( .A0(\memory[21][60] ), .A1(out_new[60]), .S(N4101), .Z(n821)
         );
  CMX2X4 U3897 ( .A0(\memory[21][59] ), .A1(out_new[59]), .S(N4101), .Z(n822)
         );
  CMX2X4 U3898 ( .A0(\memory[21][58] ), .A1(out_new[58]), .S(N4101), .Z(n823)
         );
  CMX2X4 U3899 ( .A0(\memory[21][57] ), .A1(out_new[57]), .S(N4101), .Z(n824)
         );
  CMX2X4 U3900 ( .A0(\memory[21][56] ), .A1(out_new[56]), .S(N4101), .Z(n825)
         );
  CMX2X4 U3901 ( .A0(\memory[21][55] ), .A1(out_new[55]), .S(N4101), .Z(n826)
         );
  CMX2X4 U3902 ( .A0(\memory[21][54] ), .A1(out_new[54]), .S(N4101), .Z(n827)
         );
  CMX2X4 U3903 ( .A0(\memory[21][53] ), .A1(out_new[53]), .S(N4101), .Z(n828)
         );
  CMX2X4 U3904 ( .A0(\memory[21][52] ), .A1(out_new[52]), .S(N4101), .Z(n829)
         );
  CMX2X4 U3905 ( .A0(\memory[21][51] ), .A1(out_new[51]), .S(N4101), .Z(n830)
         );
  CMX2X4 U3906 ( .A0(\memory[21][50] ), .A1(out_new[50]), .S(N4101), .Z(n831)
         );
  CMX2X4 U3907 ( .A0(\memory[21][49] ), .A1(out_new[49]), .S(N4101), .Z(n832)
         );
  CMX2X4 U3908 ( .A0(\memory[21][48] ), .A1(out_new[48]), .S(N4101), .Z(n833)
         );
  CMX2X4 U3909 ( .A0(\memory[21][47] ), .A1(out_new[47]), .S(N4101), .Z(n834)
         );
  CMX2X4 U3910 ( .A0(\memory[21][46] ), .A1(out_new[46]), .S(N4101), .Z(n835)
         );
  CMX2X4 U3911 ( .A0(\memory[21][45] ), .A1(out_new[45]), .S(N4101), .Z(n836)
         );
  CMX2X4 U3912 ( .A0(\memory[21][44] ), .A1(out_new[44]), .S(N4101), .Z(n837)
         );
  CMX2X4 U3913 ( .A0(\memory[21][43] ), .A1(out_new[43]), .S(N4101), .Z(n838)
         );
  CMX2X4 U3914 ( .A0(\memory[21][42] ), .A1(out_new[42]), .S(N4101), .Z(n839)
         );
  CMX2X4 U3915 ( .A0(\memory[21][41] ), .A1(out_new[41]), .S(N4101), .Z(n840)
         );
  CMX2X4 U3916 ( .A0(\memory[21][40] ), .A1(out_new[40]), .S(N4101), .Z(n841)
         );
  CMX2X4 U3917 ( .A0(\memory[21][39] ), .A1(out_new[39]), .S(N4101), .Z(n842)
         );
  CMX2X4 U3918 ( .A0(\memory[21][38] ), .A1(out_new[38]), .S(N4101), .Z(n843)
         );
  CMX2X4 U3919 ( .A0(\memory[21][37] ), .A1(out_new[37]), .S(N4101), .Z(n844)
         );
  CMX2X4 U3920 ( .A0(\memory[21][36] ), .A1(out_new[36]), .S(N4101), .Z(n845)
         );
  CMX2X4 U3921 ( .A0(\memory[21][35] ), .A1(out_new[35]), .S(N4101), .Z(n846)
         );
  CMX2X4 U3922 ( .A0(\memory[21][34] ), .A1(out_new[34]), .S(N4101), .Z(n847)
         );
  CMX2X4 U3923 ( .A0(\memory[21][33] ), .A1(out_new[33]), .S(N4101), .Z(n848)
         );
  CMX2X4 U3924 ( .A0(\memory[21][32] ), .A1(out_new[32]), .S(N4101), .Z(n849)
         );
  CMX2X4 U3925 ( .A0(\memory[21][31] ), .A1(out_new[31]), .S(N4101), .Z(n850)
         );
  CMX2X4 U3926 ( .A0(\memory[21][30] ), .A1(out_new[30]), .S(N4101), .Z(n851)
         );
  CMX2X4 U3927 ( .A0(\memory[21][29] ), .A1(out_new[29]), .S(N4101), .Z(n852)
         );
  CMX2X4 U3928 ( .A0(\memory[21][28] ), .A1(out_new[28]), .S(N4101), .Z(n853)
         );
  CMX2X4 U3929 ( .A0(\memory[21][27] ), .A1(out_new[27]), .S(N4101), .Z(n854)
         );
  CMX2X4 U3930 ( .A0(\memory[21][26] ), .A1(out_new[26]), .S(N4101), .Z(n855)
         );
  CMX2X4 U3931 ( .A0(\memory[21][25] ), .A1(out_new[25]), .S(N4101), .Z(n856)
         );
  CMX2X4 U3932 ( .A0(\memory[21][24] ), .A1(out_new[24]), .S(N4101), .Z(n857)
         );
  CMX2X4 U3933 ( .A0(\memory[21][23] ), .A1(out_new[23]), .S(N4101), .Z(n858)
         );
  CMX2X4 U3934 ( .A0(\memory[21][22] ), .A1(out_new[22]), .S(N4101), .Z(n859)
         );
  CMX2X4 U3935 ( .A0(\memory[21][21] ), .A1(out_new[21]), .S(N4101), .Z(n860)
         );
  CMX2X4 U3936 ( .A0(\memory[21][20] ), .A1(out_new[20]), .S(N4101), .Z(n861)
         );
  CMX2X4 U3937 ( .A0(\memory[21][19] ), .A1(out_new[19]), .S(N4101), .Z(n862)
         );
  CMX2X4 U3938 ( .A0(\memory[21][18] ), .A1(out_new[18]), .S(N4101), .Z(n863)
         );
  CMX2X4 U3939 ( .A0(\memory[21][17] ), .A1(out_new[17]), .S(N4101), .Z(n864)
         );
  CMX2X4 U3940 ( .A0(\memory[21][16] ), .A1(out_new[16]), .S(N4101), .Z(n865)
         );
  CMX2X4 U3941 ( .A0(\memory[21][15] ), .A1(out_new[15]), .S(N4101), .Z(n866)
         );
  CMX2X4 U3942 ( .A0(\memory[21][14] ), .A1(out_new[14]), .S(N4101), .Z(n867)
         );
  CMX2X4 U3943 ( .A0(\memory[21][13] ), .A1(out_new[13]), .S(N4101), .Z(n868)
         );
  CMX2X4 U3944 ( .A0(\memory[21][12] ), .A1(out_new[12]), .S(N4101), .Z(n869)
         );
  CMX2X4 U3945 ( .A0(\memory[21][11] ), .A1(out_new[11]), .S(N4101), .Z(n870)
         );
  CMX2X4 U3946 ( .A0(\memory[21][10] ), .A1(out_new[10]), .S(N4101), .Z(n871)
         );
  CMX2X4 U3947 ( .A0(\memory[21][9] ), .A1(out_new[9]), .S(N4101), .Z(n872) );
  CMX2X4 U3948 ( .A0(\memory[21][8] ), .A1(out_new[8]), .S(N4101), .Z(n873) );
  CMX2X4 U3949 ( .A0(\memory[21][7] ), .A1(out_new[7]), .S(N4101), .Z(n874) );
  CMX2X4 U3950 ( .A0(\memory[21][6] ), .A1(out_new[6]), .S(N4101), .Z(n875) );
  CMX2X4 U3951 ( .A0(\memory[21][5] ), .A1(out_new[5]), .S(N4101), .Z(n876) );
  CMX2X4 U3952 ( .A0(\memory[21][4] ), .A1(out_new[4]), .S(N4101), .Z(n877) );
  CMX2X4 U3953 ( .A0(\memory[21][3] ), .A1(out_new[3]), .S(N4101), .Z(n878) );
  CMX2X4 U3954 ( .A0(\memory[21][2] ), .A1(out_new[2]), .S(N4101), .Z(n879) );
  CMX2X4 U3955 ( .A0(\memory[21][1] ), .A1(out_new[1]), .S(N4101), .Z(n880) );
  CMX2X4 U3956 ( .A0(\memory[21][0] ), .A1(out_new[0]), .S(N4101), .Z(n881) );
  CMX2X2 U3957 ( .A0(\memory[20][63] ), .A1(out_new[63]), .S(N4030), .Z(n889)
         );
  CMX2X2 U3958 ( .A0(\memory[20][62] ), .A1(out_new[62]), .S(N4030), .Z(n890)
         );
  CMX2X2 U3959 ( .A0(\memory[20][61] ), .A1(out_new[61]), .S(N4030), .Z(n891)
         );
  CMX2X2 U3960 ( .A0(\memory[20][60] ), .A1(out_new[60]), .S(N4030), .Z(n892)
         );
  CMX2X2 U3961 ( .A0(\memory[20][59] ), .A1(out_new[59]), .S(N4030), .Z(n893)
         );
  CMX2X2 U3962 ( .A0(\memory[20][58] ), .A1(out_new[58]), .S(N4030), .Z(n894)
         );
  CMX2X2 U3963 ( .A0(\memory[20][57] ), .A1(out_new[57]), .S(N4030), .Z(n895)
         );
  CMX2X2 U3964 ( .A0(\memory[20][56] ), .A1(out_new[56]), .S(N4030), .Z(n896)
         );
  CMX2X2 U3965 ( .A0(\memory[20][55] ), .A1(out_new[55]), .S(N4030), .Z(n897)
         );
  CMX2X2 U3966 ( .A0(\memory[20][54] ), .A1(out_new[54]), .S(N4030), .Z(n898)
         );
  CMX2X2 U3967 ( .A0(\memory[20][53] ), .A1(out_new[53]), .S(N4030), .Z(n899)
         );
  CMX2X2 U3968 ( .A0(\memory[20][52] ), .A1(out_new[52]), .S(N4030), .Z(n900)
         );
  CMX2X2 U3969 ( .A0(\memory[20][51] ), .A1(out_new[51]), .S(N4030), .Z(n901)
         );
  CMX2X2 U3970 ( .A0(\memory[20][50] ), .A1(out_new[50]), .S(N4030), .Z(n902)
         );
  CMX2X2 U3971 ( .A0(\memory[20][49] ), .A1(out_new[49]), .S(N4030), .Z(n903)
         );
  CMX2X2 U3972 ( .A0(\memory[20][48] ), .A1(out_new[48]), .S(N4030), .Z(n904)
         );
  CMX2X2 U3973 ( .A0(\memory[20][47] ), .A1(out_new[47]), .S(N4030), .Z(n905)
         );
  CMX2X2 U3974 ( .A0(\memory[20][46] ), .A1(out_new[46]), .S(N4030), .Z(n906)
         );
  CMX2X2 U3975 ( .A0(\memory[20][45] ), .A1(out_new[45]), .S(N4030), .Z(n907)
         );
  CMX2X2 U3976 ( .A0(\memory[20][44] ), .A1(out_new[44]), .S(N4030), .Z(n908)
         );
  CMX2X2 U3977 ( .A0(\memory[20][43] ), .A1(out_new[43]), .S(N4030), .Z(n909)
         );
  CMX2X2 U3978 ( .A0(\memory[20][42] ), .A1(out_new[42]), .S(N4030), .Z(n910)
         );
  CMX2X2 U3979 ( .A0(\memory[20][41] ), .A1(out_new[41]), .S(N4030), .Z(n911)
         );
  CMX2X2 U3980 ( .A0(\memory[20][40] ), .A1(out_new[40]), .S(N4030), .Z(n912)
         );
  CMX2X2 U3981 ( .A0(\memory[20][39] ), .A1(out_new[39]), .S(N4030), .Z(n913)
         );
  CMX2X2 U3982 ( .A0(\memory[20][38] ), .A1(out_new[38]), .S(N4030), .Z(n914)
         );
  CMX2X2 U3983 ( .A0(\memory[20][37] ), .A1(out_new[37]), .S(N4030), .Z(n915)
         );
  CMX2X2 U3984 ( .A0(\memory[20][36] ), .A1(out_new[36]), .S(N4030), .Z(n916)
         );
  CMX2X2 U3985 ( .A0(\memory[20][35] ), .A1(out_new[35]), .S(N4030), .Z(n917)
         );
  CMX2X2 U3986 ( .A0(\memory[20][34] ), .A1(out_new[34]), .S(N4030), .Z(n918)
         );
  CMX2X2 U3987 ( .A0(\memory[20][33] ), .A1(out_new[33]), .S(N4030), .Z(n919)
         );
  CMX2X2 U3988 ( .A0(\memory[20][32] ), .A1(out_new[32]), .S(N4030), .Z(n920)
         );
  CMX2X2 U3989 ( .A0(\memory[20][31] ), .A1(out_new[31]), .S(N4030), .Z(n921)
         );
  CMX2X2 U3990 ( .A0(\memory[20][30] ), .A1(out_new[30]), .S(N4030), .Z(n922)
         );
  CMX2X2 U3991 ( .A0(\memory[20][29] ), .A1(out_new[29]), .S(N4030), .Z(n923)
         );
  CMX2X2 U3992 ( .A0(\memory[20][28] ), .A1(out_new[28]), .S(N4030), .Z(n924)
         );
  CMX2X2 U3993 ( .A0(\memory[20][27] ), .A1(out_new[27]), .S(N4030), .Z(n925)
         );
  CMX2X2 U3994 ( .A0(\memory[20][26] ), .A1(out_new[26]), .S(N4030), .Z(n926)
         );
  CMX2X2 U3995 ( .A0(\memory[20][25] ), .A1(out_new[25]), .S(N4030), .Z(n927)
         );
  CMX2X2 U3996 ( .A0(\memory[20][24] ), .A1(out_new[24]), .S(N4030), .Z(n928)
         );
  CMX2X2 U3997 ( .A0(\memory[20][23] ), .A1(out_new[23]), .S(N4030), .Z(n929)
         );
  CMX2X2 U3998 ( .A0(\memory[20][22] ), .A1(out_new[22]), .S(N4030), .Z(n930)
         );
  CMX2X2 U3999 ( .A0(\memory[20][21] ), .A1(out_new[21]), .S(N4030), .Z(n931)
         );
  CMX2X2 U4000 ( .A0(\memory[20][20] ), .A1(out_new[20]), .S(N4030), .Z(n932)
         );
  CMX2X2 U4001 ( .A0(\memory[20][19] ), .A1(out_new[19]), .S(N4030), .Z(n933)
         );
  CMX2X2 U4002 ( .A0(\memory[20][18] ), .A1(out_new[18]), .S(N4030), .Z(n934)
         );
  CMX2X2 U4003 ( .A0(\memory[20][17] ), .A1(out_new[17]), .S(N4030), .Z(n935)
         );
  CMX2X2 U4004 ( .A0(\memory[20][16] ), .A1(out_new[16]), .S(N4030), .Z(n936)
         );
  CMX2X2 U4005 ( .A0(\memory[20][15] ), .A1(out_new[15]), .S(N4030), .Z(n937)
         );
  CMX2X2 U4006 ( .A0(\memory[20][14] ), .A1(out_new[14]), .S(N4030), .Z(n938)
         );
  CMX2X2 U4007 ( .A0(\memory[20][13] ), .A1(out_new[13]), .S(N4030), .Z(n939)
         );
  CMX2X2 U4008 ( .A0(\memory[20][12] ), .A1(out_new[12]), .S(N4030), .Z(n940)
         );
  CMX2X2 U4009 ( .A0(\memory[20][11] ), .A1(out_new[11]), .S(N4030), .Z(n941)
         );
  CMX2X2 U4010 ( .A0(\memory[20][10] ), .A1(out_new[10]), .S(N4030), .Z(n942)
         );
  CMX2X2 U4011 ( .A0(\memory[20][9] ), .A1(out_new[9]), .S(N4030), .Z(n943) );
  CMX2X2 U4012 ( .A0(\memory[20][8] ), .A1(out_new[8]), .S(N4030), .Z(n944) );
  CMX2X2 U4013 ( .A0(\memory[20][7] ), .A1(out_new[7]), .S(N4030), .Z(n945) );
  CMX2X2 U4014 ( .A0(\memory[20][6] ), .A1(out_new[6]), .S(N4030), .Z(n946) );
  CMX2X2 U4015 ( .A0(\memory[20][5] ), .A1(out_new[5]), .S(N4030), .Z(n947) );
  CMX2X2 U4016 ( .A0(\memory[20][4] ), .A1(out_new[4]), .S(N4030), .Z(n948) );
  CMX2X2 U4017 ( .A0(\memory[20][3] ), .A1(out_new[3]), .S(N4030), .Z(n949) );
  CMX2X2 U4018 ( .A0(\memory[20][2] ), .A1(out_new[2]), .S(N4030), .Z(n950) );
  CMX2X2 U4019 ( .A0(\memory[20][1] ), .A1(out_new[1]), .S(N4030), .Z(n951) );
  CMX2X2 U4020 ( .A0(\memory[20][0] ), .A1(out_new[0]), .S(N4030), .Z(n952) );
  CMX2X2 U4021 ( .A0(\memory[18][63] ), .A1(out_new[63]), .S(N3888), .Z(n1031)
         );
  CMX2X2 U4022 ( .A0(\memory[18][62] ), .A1(out_new[62]), .S(N3888), .Z(n1032)
         );
  CMX2X2 U4023 ( .A0(\memory[18][61] ), .A1(out_new[61]), .S(N3888), .Z(n1033)
         );
  CMX2X2 U4024 ( .A0(\memory[18][60] ), .A1(out_new[60]), .S(N3888), .Z(n1034)
         );
  CMX2X2 U4025 ( .A0(\memory[18][59] ), .A1(out_new[59]), .S(N3888), .Z(n1035)
         );
  CMX2X2 U4026 ( .A0(\memory[18][58] ), .A1(out_new[58]), .S(N3888), .Z(n1036)
         );
  CMX2X2 U4027 ( .A0(\memory[18][57] ), .A1(out_new[57]), .S(N3888), .Z(n1037)
         );
  CMX2X2 U4028 ( .A0(\memory[18][56] ), .A1(out_new[56]), .S(N3888), .Z(n1038)
         );
  CMX2X2 U4029 ( .A0(\memory[18][55] ), .A1(out_new[55]), .S(N3888), .Z(n1039)
         );
  CMX2X2 U4030 ( .A0(\memory[18][54] ), .A1(out_new[54]), .S(N3888), .Z(n1040)
         );
  CMX2X2 U4031 ( .A0(\memory[18][53] ), .A1(out_new[53]), .S(N3888), .Z(n1041)
         );
  CMX2X2 U4032 ( .A0(\memory[18][52] ), .A1(out_new[52]), .S(N3888), .Z(n1042)
         );
  CMX2X2 U4033 ( .A0(\memory[18][51] ), .A1(out_new[51]), .S(N3888), .Z(n1043)
         );
  CMX2X2 U4034 ( .A0(\memory[18][50] ), .A1(out_new[50]), .S(N3888), .Z(n1044)
         );
  CMX2X2 U4035 ( .A0(\memory[18][49] ), .A1(out_new[49]), .S(N3888), .Z(n1045)
         );
  CMX2X2 U4036 ( .A0(\memory[18][48] ), .A1(out_new[48]), .S(N3888), .Z(n1046)
         );
  CMX2X2 U4037 ( .A0(\memory[18][47] ), .A1(out_new[47]), .S(N3888), .Z(n1047)
         );
  CMX2X2 U4038 ( .A0(\memory[18][46] ), .A1(out_new[46]), .S(N3888), .Z(n1048)
         );
  CMX2X2 U4039 ( .A0(\memory[18][45] ), .A1(out_new[45]), .S(N3888), .Z(n1049)
         );
  CMX2X2 U4040 ( .A0(\memory[18][44] ), .A1(out_new[44]), .S(N3888), .Z(n1050)
         );
  CMX2X2 U4041 ( .A0(\memory[18][43] ), .A1(out_new[43]), .S(N3888), .Z(n1051)
         );
  CMX2X2 U4042 ( .A0(\memory[18][42] ), .A1(out_new[42]), .S(N3888), .Z(n1052)
         );
  CMX2X2 U4043 ( .A0(\memory[18][41] ), .A1(out_new[41]), .S(N3888), .Z(n1053)
         );
  CMX2X2 U4044 ( .A0(\memory[18][40] ), .A1(out_new[40]), .S(N3888), .Z(n1054)
         );
  CMX2X2 U4045 ( .A0(\memory[18][39] ), .A1(out_new[39]), .S(N3888), .Z(n1055)
         );
  CMX2X2 U4046 ( .A0(\memory[18][38] ), .A1(out_new[38]), .S(N3888), .Z(n1056)
         );
  CMX2X2 U4047 ( .A0(\memory[18][37] ), .A1(out_new[37]), .S(N3888), .Z(n1057)
         );
  CMX2X2 U4048 ( .A0(\memory[18][36] ), .A1(out_new[36]), .S(N3888), .Z(n1058)
         );
  CMX2X2 U4049 ( .A0(\memory[18][35] ), .A1(out_new[35]), .S(N3888), .Z(n1059)
         );
  CMX2X2 U4050 ( .A0(\memory[18][34] ), .A1(out_new[34]), .S(N3888), .Z(n1060)
         );
  CMX2X2 U4051 ( .A0(\memory[18][33] ), .A1(out_new[33]), .S(N3888), .Z(n1061)
         );
  CMX2X2 U4052 ( .A0(\memory[18][32] ), .A1(out_new[32]), .S(N3888), .Z(n1062)
         );
  CMX2X2 U4053 ( .A0(\memory[18][31] ), .A1(out_new[31]), .S(N3888), .Z(n1063)
         );
  CMX2X2 U4054 ( .A0(\memory[18][30] ), .A1(out_new[30]), .S(N3888), .Z(n1064)
         );
  CMX2X2 U4055 ( .A0(\memory[18][29] ), .A1(out_new[29]), .S(N3888), .Z(n1065)
         );
  CMX2X2 U4056 ( .A0(\memory[18][28] ), .A1(out_new[28]), .S(N3888), .Z(n1066)
         );
  CMX2X2 U4057 ( .A0(\memory[18][27] ), .A1(out_new[27]), .S(N3888), .Z(n1067)
         );
  CMX2X2 U4058 ( .A0(\memory[18][26] ), .A1(out_new[26]), .S(N3888), .Z(n1068)
         );
  CMX2X2 U4059 ( .A0(\memory[18][25] ), .A1(out_new[25]), .S(N3888), .Z(n1069)
         );
  CMX2X2 U4060 ( .A0(\memory[18][24] ), .A1(out_new[24]), .S(N3888), .Z(n1070)
         );
  CMX2X2 U4061 ( .A0(\memory[18][23] ), .A1(out_new[23]), .S(N3888), .Z(n1071)
         );
  CMX2X2 U4062 ( .A0(\memory[18][22] ), .A1(out_new[22]), .S(N3888), .Z(n1072)
         );
  CMX2X2 U4063 ( .A0(\memory[18][21] ), .A1(out_new[21]), .S(N3888), .Z(n1073)
         );
  CMX2X2 U4064 ( .A0(\memory[18][20] ), .A1(out_new[20]), .S(N3888), .Z(n1074)
         );
  CMX2X2 U4065 ( .A0(\memory[18][19] ), .A1(out_new[19]), .S(N3888), .Z(n1075)
         );
  CMX2X2 U4066 ( .A0(\memory[18][18] ), .A1(out_new[18]), .S(N3888), .Z(n1076)
         );
  CMX2X2 U4067 ( .A0(\memory[18][17] ), .A1(out_new[17]), .S(N3888), .Z(n1077)
         );
  CMX2X2 U4068 ( .A0(\memory[18][16] ), .A1(out_new[16]), .S(N3888), .Z(n1078)
         );
  CMX2X2 U4069 ( .A0(\memory[18][15] ), .A1(out_new[15]), .S(N3888), .Z(n1079)
         );
  CMX2X2 U4070 ( .A0(\memory[18][14] ), .A1(out_new[14]), .S(N3888), .Z(n1080)
         );
  CMX2X2 U4071 ( .A0(\memory[18][13] ), .A1(out_new[13]), .S(N3888), .Z(n1081)
         );
  CMX2X2 U4072 ( .A0(\memory[18][12] ), .A1(out_new[12]), .S(N3888), .Z(n1082)
         );
  CMX2X2 U4073 ( .A0(\memory[18][11] ), .A1(out_new[11]), .S(N3888), .Z(n1083)
         );
  CMX2X2 U4074 ( .A0(\memory[18][10] ), .A1(out_new[10]), .S(N3888), .Z(n1084)
         );
  CMX2X2 U4075 ( .A0(\memory[18][9] ), .A1(out_new[9]), .S(N3888), .Z(n1085)
         );
  CMX2X2 U4076 ( .A0(\memory[18][8] ), .A1(out_new[8]), .S(N3888), .Z(n1086)
         );
  CMX2X2 U4077 ( .A0(\memory[18][7] ), .A1(out_new[7]), .S(N3888), .Z(n1087)
         );
  CMX2X2 U4078 ( .A0(\memory[18][6] ), .A1(out_new[6]), .S(N3888), .Z(n1088)
         );
  CMX2X2 U4079 ( .A0(\memory[18][5] ), .A1(out_new[5]), .S(N3888), .Z(n1089)
         );
  CMX2X2 U4080 ( .A0(\memory[18][4] ), .A1(out_new[4]), .S(N3888), .Z(n1090)
         );
  CMX2X2 U4081 ( .A0(\memory[18][3] ), .A1(out_new[3]), .S(N3888), .Z(n1091)
         );
  CMX2X2 U4082 ( .A0(\memory[18][2] ), .A1(out_new[2]), .S(N3888), .Z(n1092)
         );
  CMX2X2 U4083 ( .A0(\memory[18][1] ), .A1(out_new[1]), .S(N3888), .Z(n1093)
         );
  CMX2X2 U4084 ( .A0(\memory[18][0] ), .A1(out_new[0]), .S(N3888), .Z(n1094)
         );
  CMX2X2 U4085 ( .A0(\memory[17][63] ), .A1(out_new[63]), .S(N3817), .Z(n1102)
         );
  CMX2X2 U4086 ( .A0(\memory[17][62] ), .A1(out_new[62]), .S(N3817), .Z(n1103)
         );
  CMX2X2 U4087 ( .A0(\memory[17][61] ), .A1(out_new[61]), .S(N3817), .Z(n1104)
         );
  CMX2X2 U4088 ( .A0(\memory[17][60] ), .A1(out_new[60]), .S(N3817), .Z(n1105)
         );
  CMX2X2 U4089 ( .A0(\memory[17][59] ), .A1(out_new[59]), .S(N3817), .Z(n1106)
         );
  CMX2X2 U4090 ( .A0(\memory[17][58] ), .A1(out_new[58]), .S(N3817), .Z(n1107)
         );
  CMX2X2 U4091 ( .A0(\memory[17][57] ), .A1(out_new[57]), .S(N3817), .Z(n1108)
         );
  CMX2X2 U4092 ( .A0(\memory[17][56] ), .A1(out_new[56]), .S(N3817), .Z(n1109)
         );
  CMX2X2 U4093 ( .A0(\memory[17][55] ), .A1(out_new[55]), .S(N3817), .Z(n1110)
         );
  CMX2X2 U4094 ( .A0(\memory[17][54] ), .A1(out_new[54]), .S(N3817), .Z(n1111)
         );
  CMX2X2 U4095 ( .A0(\memory[17][53] ), .A1(out_new[53]), .S(N3817), .Z(n1112)
         );
  CMX2X2 U4096 ( .A0(\memory[17][52] ), .A1(out_new[52]), .S(N3817), .Z(n1113)
         );
  CMX2X2 U4097 ( .A0(\memory[17][51] ), .A1(out_new[51]), .S(N3817), .Z(n1114)
         );
  CMX2X2 U4098 ( .A0(\memory[17][50] ), .A1(out_new[50]), .S(N3817), .Z(n1115)
         );
  CMX2X2 U4099 ( .A0(\memory[17][49] ), .A1(out_new[49]), .S(N3817), .Z(n1116)
         );
  CMX2X2 U4100 ( .A0(\memory[17][48] ), .A1(out_new[48]), .S(N3817), .Z(n1117)
         );
  CMX2X2 U4101 ( .A0(\memory[17][47] ), .A1(out_new[47]), .S(N3817), .Z(n1118)
         );
  CMX2X2 U4102 ( .A0(\memory[17][46] ), .A1(out_new[46]), .S(N3817), .Z(n1119)
         );
  CMX2X2 U4103 ( .A0(\memory[17][45] ), .A1(out_new[45]), .S(N3817), .Z(n1120)
         );
  CMX2X2 U4104 ( .A0(\memory[17][44] ), .A1(out_new[44]), .S(N3817), .Z(n1121)
         );
  CMX2X2 U4105 ( .A0(\memory[17][43] ), .A1(out_new[43]), .S(N3817), .Z(n1122)
         );
  CMX2X2 U4106 ( .A0(\memory[17][42] ), .A1(out_new[42]), .S(N3817), .Z(n1123)
         );
  CMX2X2 U4107 ( .A0(\memory[17][41] ), .A1(out_new[41]), .S(N3817), .Z(n1124)
         );
  CMX2X2 U4108 ( .A0(\memory[17][40] ), .A1(out_new[40]), .S(N3817), .Z(n1125)
         );
  CMX2X2 U4109 ( .A0(\memory[17][39] ), .A1(out_new[39]), .S(N3817), .Z(n1126)
         );
  CMX2X2 U4110 ( .A0(\memory[17][38] ), .A1(out_new[38]), .S(N3817), .Z(n1127)
         );
  CMX2X2 U4111 ( .A0(\memory[17][37] ), .A1(out_new[37]), .S(N3817), .Z(n1128)
         );
  CMX2X2 U4112 ( .A0(\memory[17][36] ), .A1(out_new[36]), .S(N3817), .Z(n1129)
         );
  CMX2X2 U4113 ( .A0(\memory[17][35] ), .A1(out_new[35]), .S(N3817), .Z(n1130)
         );
  CMX2X2 U4114 ( .A0(\memory[17][34] ), .A1(out_new[34]), .S(N3817), .Z(n1131)
         );
  CMX2X2 U4115 ( .A0(\memory[17][33] ), .A1(out_new[33]), .S(N3817), .Z(n1132)
         );
  CMX2X2 U4116 ( .A0(\memory[17][32] ), .A1(out_new[32]), .S(N3817), .Z(n1133)
         );
  CMX2X2 U4117 ( .A0(\memory[17][31] ), .A1(out_new[31]), .S(N3817), .Z(n1134)
         );
  CMX2X2 U4118 ( .A0(\memory[17][30] ), .A1(out_new[30]), .S(N3817), .Z(n1135)
         );
  CMX2X2 U4119 ( .A0(\memory[17][29] ), .A1(out_new[29]), .S(N3817), .Z(n1136)
         );
  CMX2X2 U4120 ( .A0(\memory[17][28] ), .A1(out_new[28]), .S(N3817), .Z(n1137)
         );
  CMX2X2 U4121 ( .A0(\memory[17][27] ), .A1(out_new[27]), .S(N3817), .Z(n1138)
         );
  CMX2X2 U4122 ( .A0(\memory[17][26] ), .A1(out_new[26]), .S(N3817), .Z(n1139)
         );
  CMX2X2 U4123 ( .A0(\memory[17][25] ), .A1(out_new[25]), .S(N3817), .Z(n1140)
         );
  CMX2X2 U4124 ( .A0(\memory[17][24] ), .A1(out_new[24]), .S(N3817), .Z(n1141)
         );
  CMX2X2 U4125 ( .A0(\memory[17][23] ), .A1(out_new[23]), .S(N3817), .Z(n1142)
         );
  CMX2X2 U4126 ( .A0(\memory[17][22] ), .A1(out_new[22]), .S(N3817), .Z(n1143)
         );
  CMX2X2 U4127 ( .A0(\memory[17][21] ), .A1(out_new[21]), .S(N3817), .Z(n1144)
         );
  CMX2X2 U4128 ( .A0(\memory[17][20] ), .A1(out_new[20]), .S(N3817), .Z(n1145)
         );
  CMX2X2 U4129 ( .A0(\memory[17][19] ), .A1(out_new[19]), .S(N3817), .Z(n1146)
         );
  CMX2X2 U4130 ( .A0(\memory[17][18] ), .A1(out_new[18]), .S(N3817), .Z(n1147)
         );
  CMX2X2 U4131 ( .A0(\memory[17][17] ), .A1(out_new[17]), .S(N3817), .Z(n1148)
         );
  CMX2X2 U4132 ( .A0(\memory[17][16] ), .A1(out_new[16]), .S(N3817), .Z(n1149)
         );
  CMX2X2 U4133 ( .A0(\memory[17][15] ), .A1(out_new[15]), .S(N3817), .Z(n1150)
         );
  CMX2X2 U4134 ( .A0(\memory[17][14] ), .A1(out_new[14]), .S(N3817), .Z(n1151)
         );
  CMX2X2 U4135 ( .A0(\memory[17][13] ), .A1(out_new[13]), .S(N3817), .Z(n1152)
         );
  CMX2X2 U4136 ( .A0(\memory[17][12] ), .A1(out_new[12]), .S(N3817), .Z(n1153)
         );
  CMX2X2 U4137 ( .A0(\memory[17][11] ), .A1(out_new[11]), .S(N3817), .Z(n1154)
         );
  CMX2X2 U4138 ( .A0(\memory[17][10] ), .A1(out_new[10]), .S(N3817), .Z(n1155)
         );
  CMX2X2 U4139 ( .A0(\memory[17][9] ), .A1(out_new[9]), .S(N3817), .Z(n1156)
         );
  CMX2X2 U4140 ( .A0(\memory[17][8] ), .A1(out_new[8]), .S(N3817), .Z(n1157)
         );
  CMX2X2 U4141 ( .A0(\memory[17][7] ), .A1(out_new[7]), .S(N3817), .Z(n1158)
         );
  CMX2X2 U4142 ( .A0(\memory[17][6] ), .A1(out_new[6]), .S(N3817), .Z(n1159)
         );
  CMX2X2 U4143 ( .A0(\memory[17][5] ), .A1(out_new[5]), .S(N3817), .Z(n1160)
         );
  CMX2X2 U4144 ( .A0(\memory[17][4] ), .A1(out_new[4]), .S(N3817), .Z(n1161)
         );
  CMX2X2 U4145 ( .A0(\memory[17][3] ), .A1(out_new[3]), .S(N3817), .Z(n1162)
         );
  CMX2X2 U4146 ( .A0(\memory[17][2] ), .A1(out_new[2]), .S(N3817), .Z(n1163)
         );
  CMX2X2 U4147 ( .A0(\memory[17][1] ), .A1(out_new[1]), .S(N3817), .Z(n1164)
         );
  CMX2X2 U4148 ( .A0(\memory[17][0] ), .A1(out_new[0]), .S(N3817), .Z(n1165)
         );
  CMX2X2 U4149 ( .A0(\memory[16][63] ), .A1(out_new[63]), .S(N3746), .Z(n1173)
         );
  CMX2X2 U4150 ( .A0(\memory[16][62] ), .A1(out_new[62]), .S(N3746), .Z(n1174)
         );
  CMX2X2 U4151 ( .A0(\memory[16][61] ), .A1(out_new[61]), .S(N3746), .Z(n1175)
         );
  CMX2X2 U4152 ( .A0(\memory[16][60] ), .A1(out_new[60]), .S(N3746), .Z(n1176)
         );
  CMX2X2 U4153 ( .A0(\memory[16][59] ), .A1(out_new[59]), .S(N3746), .Z(n1177)
         );
  CMX2X2 U4154 ( .A0(\memory[16][58] ), .A1(out_new[58]), .S(N3746), .Z(n1178)
         );
  CMX2X2 U4155 ( .A0(\memory[16][57] ), .A1(out_new[57]), .S(N3746), .Z(n1179)
         );
  CMX2X2 U4156 ( .A0(\memory[16][56] ), .A1(out_new[56]), .S(N3746), .Z(n1180)
         );
  CMX2X2 U4157 ( .A0(\memory[16][55] ), .A1(out_new[55]), .S(N3746), .Z(n1181)
         );
  CMX2X2 U4158 ( .A0(\memory[16][54] ), .A1(out_new[54]), .S(N3746), .Z(n1182)
         );
  CMX2X2 U4159 ( .A0(\memory[16][53] ), .A1(out_new[53]), .S(N3746), .Z(n1183)
         );
  CMX2X2 U4160 ( .A0(\memory[16][52] ), .A1(out_new[52]), .S(N3746), .Z(n1184)
         );
  CMX2X2 U4161 ( .A0(\memory[16][51] ), .A1(out_new[51]), .S(N3746), .Z(n1185)
         );
  CMX2X2 U4162 ( .A0(\memory[16][50] ), .A1(out_new[50]), .S(N3746), .Z(n1186)
         );
  CMX2X2 U4163 ( .A0(\memory[16][49] ), .A1(out_new[49]), .S(N3746), .Z(n1187)
         );
  CMX2X2 U4164 ( .A0(\memory[16][48] ), .A1(out_new[48]), .S(N3746), .Z(n1188)
         );
  CMX2X2 U4165 ( .A0(\memory[16][47] ), .A1(out_new[47]), .S(N3746), .Z(n1189)
         );
  CMX2X2 U4166 ( .A0(\memory[16][46] ), .A1(out_new[46]), .S(N3746), .Z(n1190)
         );
  CMX2X2 U4167 ( .A0(\memory[16][45] ), .A1(out_new[45]), .S(N3746), .Z(n1191)
         );
  CMX2X2 U4168 ( .A0(\memory[16][44] ), .A1(out_new[44]), .S(N3746), .Z(n1192)
         );
  CMX2X2 U4169 ( .A0(\memory[16][43] ), .A1(out_new[43]), .S(N3746), .Z(n1193)
         );
  CMX2X2 U4170 ( .A0(\memory[16][42] ), .A1(out_new[42]), .S(N3746), .Z(n1194)
         );
  CMX2X2 U4171 ( .A0(\memory[16][41] ), .A1(out_new[41]), .S(N3746), .Z(n1195)
         );
  CMX2X2 U4172 ( .A0(\memory[16][40] ), .A1(out_new[40]), .S(N3746), .Z(n1196)
         );
  CMX2X2 U4173 ( .A0(\memory[16][39] ), .A1(out_new[39]), .S(N3746), .Z(n1197)
         );
  CMX2X2 U4174 ( .A0(\memory[16][38] ), .A1(out_new[38]), .S(N3746), .Z(n1198)
         );
  CMX2X2 U4175 ( .A0(\memory[16][37] ), .A1(out_new[37]), .S(N3746), .Z(n1199)
         );
  CMX2X2 U4176 ( .A0(\memory[16][36] ), .A1(out_new[36]), .S(N3746), .Z(n1200)
         );
  CMX2X2 U4177 ( .A0(\memory[16][35] ), .A1(out_new[35]), .S(N3746), .Z(n1201)
         );
  CMX2X2 U4178 ( .A0(\memory[16][34] ), .A1(out_new[34]), .S(N3746), .Z(n1202)
         );
  CMX2X2 U4179 ( .A0(\memory[16][33] ), .A1(out_new[33]), .S(N3746), .Z(n1203)
         );
  CMX2X2 U4180 ( .A0(\memory[16][32] ), .A1(out_new[32]), .S(N3746), .Z(n1204)
         );
  CMX2X2 U4181 ( .A0(\memory[16][31] ), .A1(out_new[31]), .S(N3746), .Z(n1205)
         );
  CMX2X2 U4182 ( .A0(\memory[16][30] ), .A1(out_new[30]), .S(N3746), .Z(n1206)
         );
  CMX2X2 U4183 ( .A0(\memory[16][29] ), .A1(out_new[29]), .S(N3746), .Z(n1207)
         );
  CMX2X2 U4184 ( .A0(\memory[16][28] ), .A1(out_new[28]), .S(N3746), .Z(n1208)
         );
  CMX2X2 U4185 ( .A0(\memory[16][27] ), .A1(out_new[27]), .S(N3746), .Z(n1209)
         );
  CMX2X2 U4186 ( .A0(\memory[16][26] ), .A1(out_new[26]), .S(N3746), .Z(n1210)
         );
  CMX2X2 U4187 ( .A0(\memory[16][25] ), .A1(out_new[25]), .S(N3746), .Z(n1211)
         );
  CMX2X2 U4188 ( .A0(\memory[16][24] ), .A1(out_new[24]), .S(N3746), .Z(n1212)
         );
  CMX2X2 U4189 ( .A0(\memory[16][23] ), .A1(out_new[23]), .S(N3746), .Z(n1213)
         );
  CMX2X2 U4190 ( .A0(\memory[16][22] ), .A1(out_new[22]), .S(N3746), .Z(n1214)
         );
  CMX2X2 U4191 ( .A0(\memory[16][21] ), .A1(out_new[21]), .S(N3746), .Z(n1215)
         );
  CMX2X2 U4192 ( .A0(\memory[16][20] ), .A1(out_new[20]), .S(N3746), .Z(n1216)
         );
  CMX2X2 U4193 ( .A0(\memory[16][19] ), .A1(out_new[19]), .S(N3746), .Z(n1217)
         );
  CMX2X2 U4194 ( .A0(\memory[16][18] ), .A1(out_new[18]), .S(N3746), .Z(n1218)
         );
  CMX2X2 U4195 ( .A0(\memory[16][17] ), .A1(out_new[17]), .S(N3746), .Z(n1219)
         );
  CMX2X2 U4196 ( .A0(\memory[16][16] ), .A1(out_new[16]), .S(N3746), .Z(n1220)
         );
  CMX2X2 U4197 ( .A0(\memory[16][15] ), .A1(out_new[15]), .S(N3746), .Z(n1221)
         );
  CMX2X2 U4198 ( .A0(\memory[16][14] ), .A1(out_new[14]), .S(N3746), .Z(n1222)
         );
  CMX2X2 U4199 ( .A0(\memory[16][13] ), .A1(out_new[13]), .S(N3746), .Z(n1223)
         );
  CMX2X2 U4200 ( .A0(\memory[16][12] ), .A1(out_new[12]), .S(N3746), .Z(n1224)
         );
  CMX2X2 U4201 ( .A0(\memory[16][11] ), .A1(out_new[11]), .S(N3746), .Z(n1225)
         );
  CMX2X2 U4202 ( .A0(\memory[16][10] ), .A1(out_new[10]), .S(N3746), .Z(n1226)
         );
  CMX2X2 U4203 ( .A0(\memory[16][9] ), .A1(out_new[9]), .S(N3746), .Z(n1227)
         );
  CMX2X2 U4204 ( .A0(\memory[16][8] ), .A1(out_new[8]), .S(N3746), .Z(n1228)
         );
  CMX2X2 U4205 ( .A0(\memory[16][7] ), .A1(out_new[7]), .S(N3746), .Z(n1229)
         );
  CMX2X2 U4206 ( .A0(\memory[16][6] ), .A1(out_new[6]), .S(N3746), .Z(n1230)
         );
  CMX2X2 U4207 ( .A0(\memory[16][5] ), .A1(out_new[5]), .S(N3746), .Z(n1231)
         );
  CMX2X2 U4208 ( .A0(\memory[16][4] ), .A1(out_new[4]), .S(N3746), .Z(n1232)
         );
  CMX2X2 U4209 ( .A0(\memory[16][3] ), .A1(out_new[3]), .S(N3746), .Z(n1233)
         );
  CMX2X2 U4210 ( .A0(\memory[16][2] ), .A1(out_new[2]), .S(N3746), .Z(n1234)
         );
  CMX2X2 U4211 ( .A0(\memory[16][1] ), .A1(out_new[1]), .S(N3746), .Z(n1235)
         );
  CMX2X2 U4212 ( .A0(\memory[16][0] ), .A1(out_new[0]), .S(N3746), .Z(n1236)
         );
  CMX2X2 U4213 ( .A0(\memory[14][63] ), .A1(out_new[63]), .S(N3604), .Z(n1315)
         );
  CMX2X2 U4214 ( .A0(\memory[14][62] ), .A1(out_new[62]), .S(N3604), .Z(n1316)
         );
  CMX2X2 U4215 ( .A0(\memory[14][61] ), .A1(out_new[61]), .S(N3604), .Z(n1317)
         );
  CMX2X2 U4216 ( .A0(\memory[14][60] ), .A1(out_new[60]), .S(N3604), .Z(n1318)
         );
  CMX2X2 U4217 ( .A0(\memory[14][59] ), .A1(out_new[59]), .S(N3604), .Z(n1319)
         );
  CMX2X2 U4218 ( .A0(\memory[14][58] ), .A1(out_new[58]), .S(N3604), .Z(n1320)
         );
  CMX2X2 U4219 ( .A0(\memory[14][57] ), .A1(out_new[57]), .S(N3604), .Z(n1321)
         );
  CMX2X2 U4220 ( .A0(\memory[14][56] ), .A1(out_new[56]), .S(N3604), .Z(n1322)
         );
  CMX2X2 U4221 ( .A0(\memory[14][55] ), .A1(out_new[55]), .S(N3604), .Z(n1323)
         );
  CMX2X2 U4222 ( .A0(\memory[14][54] ), .A1(out_new[54]), .S(N3604), .Z(n1324)
         );
  CMX2X2 U4223 ( .A0(\memory[14][53] ), .A1(out_new[53]), .S(N3604), .Z(n1325)
         );
  CMX2X2 U4224 ( .A0(\memory[14][52] ), .A1(out_new[52]), .S(N3604), .Z(n1326)
         );
  CMX2X2 U4225 ( .A0(\memory[14][51] ), .A1(out_new[51]), .S(N3604), .Z(n1327)
         );
  CMX2X2 U4226 ( .A0(\memory[14][50] ), .A1(out_new[50]), .S(N3604), .Z(n1328)
         );
  CMX2X2 U4227 ( .A0(\memory[14][49] ), .A1(out_new[49]), .S(N3604), .Z(n1329)
         );
  CMX2X2 U4228 ( .A0(\memory[14][48] ), .A1(out_new[48]), .S(N3604), .Z(n1330)
         );
  CMX2X2 U4229 ( .A0(\memory[14][47] ), .A1(out_new[47]), .S(N3604), .Z(n1331)
         );
  CMX2X2 U4230 ( .A0(\memory[14][46] ), .A1(out_new[46]), .S(N3604), .Z(n1332)
         );
  CMX2X2 U4231 ( .A0(\memory[14][45] ), .A1(out_new[45]), .S(N3604), .Z(n1333)
         );
  CMX2X2 U4232 ( .A0(\memory[14][44] ), .A1(out_new[44]), .S(N3604), .Z(n1334)
         );
  CMX2X2 U4233 ( .A0(\memory[14][43] ), .A1(out_new[43]), .S(N3604), .Z(n1335)
         );
  CMX2X2 U4234 ( .A0(\memory[14][42] ), .A1(out_new[42]), .S(N3604), .Z(n1336)
         );
  CMX2X2 U4235 ( .A0(\memory[14][41] ), .A1(out_new[41]), .S(N3604), .Z(n1337)
         );
  CMX2X2 U4236 ( .A0(\memory[14][40] ), .A1(out_new[40]), .S(N3604), .Z(n1338)
         );
  CMX2X2 U4237 ( .A0(\memory[14][39] ), .A1(out_new[39]), .S(N3604), .Z(n1339)
         );
  CMX2X2 U4238 ( .A0(\memory[14][38] ), .A1(out_new[38]), .S(N3604), .Z(n1340)
         );
  CMX2X2 U4239 ( .A0(\memory[14][37] ), .A1(out_new[37]), .S(N3604), .Z(n1341)
         );
  CMX2X2 U4240 ( .A0(\memory[14][36] ), .A1(out_new[36]), .S(N3604), .Z(n1342)
         );
  CMX2X2 U4241 ( .A0(\memory[14][35] ), .A1(out_new[35]), .S(N3604), .Z(n1343)
         );
  CMX2X2 U4242 ( .A0(\memory[14][34] ), .A1(out_new[34]), .S(N3604), .Z(n1344)
         );
  CMX2X2 U4243 ( .A0(\memory[14][33] ), .A1(out_new[33]), .S(N3604), .Z(n1345)
         );
  CMX2X2 U4244 ( .A0(\memory[14][32] ), .A1(out_new[32]), .S(N3604), .Z(n1346)
         );
  CMX2X2 U4245 ( .A0(\memory[14][31] ), .A1(out_new[31]), .S(N3604), .Z(n1347)
         );
  CMX2X2 U4246 ( .A0(\memory[14][30] ), .A1(out_new[30]), .S(N3604), .Z(n1348)
         );
  CMX2X2 U4247 ( .A0(\memory[14][29] ), .A1(out_new[29]), .S(N3604), .Z(n1349)
         );
  CMX2X2 U4248 ( .A0(\memory[14][28] ), .A1(out_new[28]), .S(N3604), .Z(n1350)
         );
  CMX2X2 U4249 ( .A0(\memory[14][27] ), .A1(out_new[27]), .S(N3604), .Z(n1351)
         );
  CMX2X2 U4250 ( .A0(\memory[14][26] ), .A1(out_new[26]), .S(N3604), .Z(n1352)
         );
  CMX2X2 U4251 ( .A0(\memory[14][25] ), .A1(out_new[25]), .S(N3604), .Z(n1353)
         );
  CMX2X2 U4252 ( .A0(\memory[14][24] ), .A1(out_new[24]), .S(N3604), .Z(n1354)
         );
  CMX2X2 U4253 ( .A0(\memory[14][23] ), .A1(out_new[23]), .S(N3604), .Z(n1355)
         );
  CMX2X2 U4254 ( .A0(\memory[14][22] ), .A1(out_new[22]), .S(N3604), .Z(n1356)
         );
  CMX2X2 U4255 ( .A0(\memory[14][21] ), .A1(out_new[21]), .S(N3604), .Z(n1357)
         );
  CMX2X2 U4256 ( .A0(\memory[14][20] ), .A1(out_new[20]), .S(N3604), .Z(n1358)
         );
  CMX2X2 U4257 ( .A0(\memory[14][19] ), .A1(out_new[19]), .S(N3604), .Z(n1359)
         );
  CMX2X2 U4258 ( .A0(\memory[14][18] ), .A1(out_new[18]), .S(N3604), .Z(n1360)
         );
  CMX2X2 U4259 ( .A0(\memory[14][17] ), .A1(out_new[17]), .S(N3604), .Z(n1361)
         );
  CMX2X2 U4260 ( .A0(\memory[14][16] ), .A1(out_new[16]), .S(N3604), .Z(n1362)
         );
  CMX2X2 U4261 ( .A0(\memory[14][15] ), .A1(out_new[15]), .S(N3604), .Z(n1363)
         );
  CMX2X2 U4262 ( .A0(\memory[14][14] ), .A1(out_new[14]), .S(N3604), .Z(n1364)
         );
  CMX2X2 U4263 ( .A0(\memory[14][13] ), .A1(out_new[13]), .S(N3604), .Z(n1365)
         );
  CMX2X2 U4264 ( .A0(\memory[14][12] ), .A1(out_new[12]), .S(N3604), .Z(n1366)
         );
  CMX2X2 U4265 ( .A0(\memory[14][11] ), .A1(out_new[11]), .S(N3604), .Z(n1367)
         );
  CMX2X2 U4266 ( .A0(\memory[14][10] ), .A1(out_new[10]), .S(N3604), .Z(n1368)
         );
  CMX2X2 U4267 ( .A0(\memory[14][9] ), .A1(out_new[9]), .S(N3604), .Z(n1369)
         );
  CMX2X2 U4268 ( .A0(\memory[14][8] ), .A1(out_new[8]), .S(N3604), .Z(n1370)
         );
  CMX2X2 U4269 ( .A0(\memory[14][7] ), .A1(out_new[7]), .S(N3604), .Z(n1371)
         );
  CMX2X2 U4270 ( .A0(\memory[14][6] ), .A1(out_new[6]), .S(N3604), .Z(n1372)
         );
  CMX2X2 U4271 ( .A0(\memory[14][5] ), .A1(out_new[5]), .S(N3604), .Z(n1373)
         );
  CMX2X2 U4272 ( .A0(\memory[14][4] ), .A1(out_new[4]), .S(N3604), .Z(n1374)
         );
  CMX2X2 U4273 ( .A0(\memory[14][3] ), .A1(out_new[3]), .S(N3604), .Z(n1375)
         );
  CMX2X2 U4274 ( .A0(\memory[14][2] ), .A1(out_new[2]), .S(N3604), .Z(n1376)
         );
  CMX2X2 U4275 ( .A0(\memory[14][1] ), .A1(out_new[1]), .S(N3604), .Z(n1377)
         );
  CMX2X2 U4276 ( .A0(\memory[14][0] ), .A1(out_new[0]), .S(N3604), .Z(n1378)
         );
  CMX2X4 U4277 ( .A0(\memory[13][63] ), .A1(out_new[63]), .S(N3533), .Z(n1386)
         );
  CMX2X4 U4278 ( .A0(\memory[13][62] ), .A1(out_new[62]), .S(N3533), .Z(n1387)
         );
  CMX2X4 U4279 ( .A0(\memory[13][61] ), .A1(out_new[61]), .S(N3533), .Z(n1388)
         );
  CMX2X4 U4280 ( .A0(\memory[13][60] ), .A1(out_new[60]), .S(N3533), .Z(n1389)
         );
  CMX2X4 U4281 ( .A0(\memory[13][59] ), .A1(out_new[59]), .S(N3533), .Z(n1390)
         );
  CMX2X4 U4282 ( .A0(\memory[13][58] ), .A1(out_new[58]), .S(N3533), .Z(n1391)
         );
  CMX2X4 U4283 ( .A0(\memory[13][57] ), .A1(out_new[57]), .S(N3533), .Z(n1392)
         );
  CMX2X4 U4284 ( .A0(\memory[13][56] ), .A1(out_new[56]), .S(N3533), .Z(n1393)
         );
  CMX2X4 U4285 ( .A0(\memory[13][55] ), .A1(out_new[55]), .S(N3533), .Z(n1394)
         );
  CMX2X4 U4286 ( .A0(\memory[13][54] ), .A1(out_new[54]), .S(N3533), .Z(n1395)
         );
  CMX2X4 U4287 ( .A0(\memory[13][53] ), .A1(out_new[53]), .S(N3533), .Z(n1396)
         );
  CMX2X4 U4288 ( .A0(\memory[13][52] ), .A1(out_new[52]), .S(N3533), .Z(n1397)
         );
  CMX2X4 U4289 ( .A0(\memory[13][51] ), .A1(out_new[51]), .S(N3533), .Z(n1398)
         );
  CMX2X4 U4290 ( .A0(\memory[13][50] ), .A1(out_new[50]), .S(N3533), .Z(n1399)
         );
  CMX2X4 U4291 ( .A0(\memory[13][49] ), .A1(out_new[49]), .S(N3533), .Z(n1400)
         );
  CMX2X4 U4292 ( .A0(\memory[13][48] ), .A1(out_new[48]), .S(N3533), .Z(n1401)
         );
  CMX2X4 U4293 ( .A0(\memory[13][47] ), .A1(out_new[47]), .S(N3533), .Z(n1402)
         );
  CMX2X4 U4294 ( .A0(\memory[13][46] ), .A1(out_new[46]), .S(N3533), .Z(n1403)
         );
  CMX2X4 U4295 ( .A0(\memory[13][45] ), .A1(out_new[45]), .S(N3533), .Z(n1404)
         );
  CMX2X4 U4296 ( .A0(\memory[13][44] ), .A1(out_new[44]), .S(N3533), .Z(n1405)
         );
  CMX2X4 U4297 ( .A0(\memory[13][43] ), .A1(out_new[43]), .S(N3533), .Z(n1406)
         );
  CMX2X4 U4298 ( .A0(\memory[13][42] ), .A1(out_new[42]), .S(N3533), .Z(n1407)
         );
  CMX2X4 U4299 ( .A0(\memory[13][41] ), .A1(out_new[41]), .S(N3533), .Z(n1408)
         );
  CMX2X4 U4300 ( .A0(\memory[13][40] ), .A1(out_new[40]), .S(N3533), .Z(n1409)
         );
  CMX2X4 U4301 ( .A0(\memory[13][39] ), .A1(out_new[39]), .S(N3533), .Z(n1410)
         );
  CMX2X4 U4302 ( .A0(\memory[13][38] ), .A1(out_new[38]), .S(N3533), .Z(n1411)
         );
  CMX2X4 U4303 ( .A0(\memory[13][37] ), .A1(out_new[37]), .S(N3533), .Z(n1412)
         );
  CMX2X4 U4304 ( .A0(\memory[13][36] ), .A1(out_new[36]), .S(N3533), .Z(n1413)
         );
  CMX2X4 U4305 ( .A0(\memory[13][35] ), .A1(out_new[35]), .S(N3533), .Z(n1414)
         );
  CMX2X4 U4306 ( .A0(\memory[13][34] ), .A1(out_new[34]), .S(N3533), .Z(n1415)
         );
  CMX2X4 U4307 ( .A0(\memory[13][33] ), .A1(out_new[33]), .S(N3533), .Z(n1416)
         );
  CMX2X4 U4308 ( .A0(\memory[13][32] ), .A1(out_new[32]), .S(N3533), .Z(n1417)
         );
  CMX2X4 U4309 ( .A0(\memory[13][31] ), .A1(out_new[31]), .S(N3533), .Z(n1418)
         );
  CMX2X4 U4310 ( .A0(\memory[13][30] ), .A1(out_new[30]), .S(N3533), .Z(n1419)
         );
  CMX2X4 U4311 ( .A0(\memory[13][29] ), .A1(out_new[29]), .S(N3533), .Z(n1420)
         );
  CMX2X4 U4312 ( .A0(\memory[13][28] ), .A1(out_new[28]), .S(N3533), .Z(n1421)
         );
  CMX2X4 U4313 ( .A0(\memory[13][27] ), .A1(out_new[27]), .S(N3533), .Z(n1422)
         );
  CMX2X4 U4314 ( .A0(\memory[13][26] ), .A1(out_new[26]), .S(N3533), .Z(n1423)
         );
  CMX2X4 U4315 ( .A0(\memory[13][25] ), .A1(out_new[25]), .S(N3533), .Z(n1424)
         );
  CMX2X4 U4316 ( .A0(\memory[13][24] ), .A1(out_new[24]), .S(N3533), .Z(n1425)
         );
  CMX2X4 U4317 ( .A0(\memory[13][23] ), .A1(out_new[23]), .S(N3533), .Z(n1426)
         );
  CMX2X4 U4318 ( .A0(\memory[13][22] ), .A1(out_new[22]), .S(N3533), .Z(n1427)
         );
  CMX2X4 U4319 ( .A0(\memory[13][21] ), .A1(out_new[21]), .S(N3533), .Z(n1428)
         );
  CMX2X4 U4320 ( .A0(\memory[13][20] ), .A1(out_new[20]), .S(N3533), .Z(n1429)
         );
  CMX2X4 U4321 ( .A0(\memory[13][19] ), .A1(out_new[19]), .S(N3533), .Z(n1430)
         );
  CMX2X4 U4322 ( .A0(\memory[13][18] ), .A1(out_new[18]), .S(N3533), .Z(n1431)
         );
  CMX2X4 U4323 ( .A0(\memory[13][17] ), .A1(out_new[17]), .S(N3533), .Z(n1432)
         );
  CMX2X4 U4324 ( .A0(\memory[13][16] ), .A1(out_new[16]), .S(N3533), .Z(n1433)
         );
  CMX2X4 U4325 ( .A0(\memory[13][15] ), .A1(out_new[15]), .S(N3533), .Z(n1434)
         );
  CMX2X4 U4326 ( .A0(\memory[13][14] ), .A1(out_new[14]), .S(N3533), .Z(n1435)
         );
  CMX2X4 U4327 ( .A0(\memory[13][13] ), .A1(out_new[13]), .S(N3533), .Z(n1436)
         );
  CMX2X4 U4328 ( .A0(\memory[13][12] ), .A1(out_new[12]), .S(N3533), .Z(n1437)
         );
  CMX2X4 U4329 ( .A0(\memory[13][11] ), .A1(out_new[11]), .S(N3533), .Z(n1438)
         );
  CMX2X4 U4330 ( .A0(\memory[13][10] ), .A1(out_new[10]), .S(N3533), .Z(n1439)
         );
  CMX2X4 U4331 ( .A0(\memory[13][9] ), .A1(out_new[9]), .S(N3533), .Z(n1440)
         );
  CMX2X4 U4332 ( .A0(\memory[13][8] ), .A1(out_new[8]), .S(N3533), .Z(n1441)
         );
  CMX2X4 U4333 ( .A0(\memory[13][7] ), .A1(out_new[7]), .S(N3533), .Z(n1442)
         );
  CMX2X4 U4334 ( .A0(\memory[13][6] ), .A1(out_new[6]), .S(N3533), .Z(n1443)
         );
  CMX2X4 U4335 ( .A0(\memory[13][5] ), .A1(out_new[5]), .S(N3533), .Z(n1444)
         );
  CMX2X4 U4336 ( .A0(\memory[13][4] ), .A1(out_new[4]), .S(N3533), .Z(n1445)
         );
  CMX2X4 U4337 ( .A0(\memory[13][3] ), .A1(out_new[3]), .S(N3533), .Z(n1446)
         );
  CMX2X4 U4338 ( .A0(\memory[13][2] ), .A1(out_new[2]), .S(N3533), .Z(n1447)
         );
  CMX2X4 U4339 ( .A0(\memory[13][1] ), .A1(out_new[1]), .S(N3533), .Z(n1448)
         );
  CMX2X4 U4340 ( .A0(\memory[13][0] ), .A1(out_new[0]), .S(N3533), .Z(n1449)
         );
  CMX2X2 U4341 ( .A0(\memory[12][63] ), .A1(out_new[63]), .S(N3462), .Z(n1457)
         );
  CMX2X2 U4342 ( .A0(\memory[12][62] ), .A1(out_new[62]), .S(N3462), .Z(n1458)
         );
  CMX2X2 U4343 ( .A0(\memory[12][61] ), .A1(out_new[61]), .S(N3462), .Z(n1459)
         );
  CMX2X2 U4344 ( .A0(\memory[12][60] ), .A1(out_new[60]), .S(N3462), .Z(n1460)
         );
  CMX2X2 U4345 ( .A0(\memory[12][59] ), .A1(out_new[59]), .S(N3462), .Z(n1461)
         );
  CMX2X2 U4346 ( .A0(\memory[12][58] ), .A1(out_new[58]), .S(N3462), .Z(n1462)
         );
  CMX2X2 U4347 ( .A0(\memory[12][57] ), .A1(out_new[57]), .S(N3462), .Z(n1463)
         );
  CMX2X2 U4348 ( .A0(\memory[12][56] ), .A1(out_new[56]), .S(N3462), .Z(n1464)
         );
  CMX2X2 U4349 ( .A0(\memory[12][55] ), .A1(out_new[55]), .S(N3462), .Z(n1465)
         );
  CMX2X2 U4350 ( .A0(\memory[12][54] ), .A1(out_new[54]), .S(N3462), .Z(n1466)
         );
  CMX2X2 U4351 ( .A0(\memory[12][53] ), .A1(out_new[53]), .S(N3462), .Z(n1467)
         );
  CMX2X2 U4352 ( .A0(\memory[12][52] ), .A1(out_new[52]), .S(N3462), .Z(n1468)
         );
  CMX2X2 U4353 ( .A0(\memory[12][51] ), .A1(out_new[51]), .S(N3462), .Z(n1469)
         );
  CMX2X2 U4354 ( .A0(\memory[12][50] ), .A1(out_new[50]), .S(N3462), .Z(n1470)
         );
  CMX2X2 U4355 ( .A0(\memory[12][49] ), .A1(out_new[49]), .S(N3462), .Z(n1471)
         );
  CMX2X2 U4356 ( .A0(\memory[12][48] ), .A1(out_new[48]), .S(N3462), .Z(n1472)
         );
  CMX2X2 U4357 ( .A0(\memory[12][47] ), .A1(out_new[47]), .S(N3462), .Z(n1473)
         );
  CMX2X2 U4358 ( .A0(\memory[12][46] ), .A1(out_new[46]), .S(N3462), .Z(n1474)
         );
  CMX2X2 U4359 ( .A0(\memory[12][45] ), .A1(out_new[45]), .S(N3462), .Z(n1475)
         );
  CMX2X2 U4360 ( .A0(\memory[12][44] ), .A1(out_new[44]), .S(N3462), .Z(n1476)
         );
  CMX2X2 U4361 ( .A0(\memory[12][43] ), .A1(out_new[43]), .S(N3462), .Z(n1477)
         );
  CMX2X2 U4362 ( .A0(\memory[12][42] ), .A1(out_new[42]), .S(N3462), .Z(n1478)
         );
  CMX2X2 U4363 ( .A0(\memory[12][41] ), .A1(out_new[41]), .S(N3462), .Z(n1479)
         );
  CMX2X2 U4364 ( .A0(\memory[12][40] ), .A1(out_new[40]), .S(N3462), .Z(n1480)
         );
  CMX2X2 U4365 ( .A0(\memory[12][39] ), .A1(out_new[39]), .S(N3462), .Z(n1481)
         );
  CMX2X2 U4366 ( .A0(\memory[12][38] ), .A1(out_new[38]), .S(N3462), .Z(n1482)
         );
  CMX2X2 U4367 ( .A0(\memory[12][37] ), .A1(out_new[37]), .S(N3462), .Z(n1483)
         );
  CMX2X2 U4368 ( .A0(\memory[12][36] ), .A1(out_new[36]), .S(N3462), .Z(n1484)
         );
  CMX2X2 U4369 ( .A0(\memory[12][35] ), .A1(out_new[35]), .S(N3462), .Z(n1485)
         );
  CMX2X2 U4370 ( .A0(\memory[12][34] ), .A1(out_new[34]), .S(N3462), .Z(n1486)
         );
  CMX2X2 U4371 ( .A0(\memory[12][33] ), .A1(out_new[33]), .S(N3462), .Z(n1487)
         );
  CMX2X2 U4372 ( .A0(\memory[12][32] ), .A1(out_new[32]), .S(N3462), .Z(n1488)
         );
  CMX2X2 U4373 ( .A0(\memory[12][31] ), .A1(out_new[31]), .S(N3462), .Z(n1489)
         );
  CMX2X2 U4374 ( .A0(\memory[12][30] ), .A1(out_new[30]), .S(N3462), .Z(n1490)
         );
  CMX2X2 U4375 ( .A0(\memory[12][29] ), .A1(out_new[29]), .S(N3462), .Z(n1491)
         );
  CMX2X2 U4376 ( .A0(\memory[12][28] ), .A1(out_new[28]), .S(N3462), .Z(n1492)
         );
  CMX2X2 U4377 ( .A0(\memory[12][27] ), .A1(out_new[27]), .S(N3462), .Z(n1493)
         );
  CMX2X2 U4378 ( .A0(\memory[12][26] ), .A1(out_new[26]), .S(N3462), .Z(n1494)
         );
  CMX2X2 U4379 ( .A0(\memory[12][25] ), .A1(out_new[25]), .S(N3462), .Z(n1495)
         );
  CMX2X2 U4380 ( .A0(\memory[12][24] ), .A1(out_new[24]), .S(N3462), .Z(n1496)
         );
  CMX2X2 U4381 ( .A0(\memory[12][23] ), .A1(out_new[23]), .S(N3462), .Z(n1497)
         );
  CMX2X2 U4382 ( .A0(\memory[12][22] ), .A1(out_new[22]), .S(N3462), .Z(n1498)
         );
  CMX2X2 U4383 ( .A0(\memory[12][21] ), .A1(out_new[21]), .S(N3462), .Z(n1499)
         );
  CMX2X2 U4384 ( .A0(\memory[12][20] ), .A1(out_new[20]), .S(N3462), .Z(n1500)
         );
  CMX2X2 U4385 ( .A0(\memory[12][19] ), .A1(out_new[19]), .S(N3462), .Z(n1501)
         );
  CMX2X2 U4386 ( .A0(\memory[12][18] ), .A1(out_new[18]), .S(N3462), .Z(n1502)
         );
  CMX2X2 U4387 ( .A0(\memory[12][17] ), .A1(out_new[17]), .S(N3462), .Z(n1503)
         );
  CMX2X2 U4388 ( .A0(\memory[12][16] ), .A1(out_new[16]), .S(N3462), .Z(n1504)
         );
  CMX2X2 U4389 ( .A0(\memory[12][15] ), .A1(out_new[15]), .S(N3462), .Z(n1505)
         );
  CMX2X2 U4390 ( .A0(\memory[12][14] ), .A1(out_new[14]), .S(N3462), .Z(n1506)
         );
  CMX2X2 U4391 ( .A0(\memory[12][13] ), .A1(out_new[13]), .S(N3462), .Z(n1507)
         );
  CMX2X2 U4392 ( .A0(\memory[12][12] ), .A1(out_new[12]), .S(N3462), .Z(n1508)
         );
  CMX2X2 U4393 ( .A0(\memory[12][11] ), .A1(out_new[11]), .S(N3462), .Z(n1509)
         );
  CMX2X2 U4394 ( .A0(\memory[12][10] ), .A1(out_new[10]), .S(N3462), .Z(n1510)
         );
  CMX2X2 U4395 ( .A0(\memory[12][9] ), .A1(out_new[9]), .S(N3462), .Z(n1511)
         );
  CMX2X2 U4396 ( .A0(\memory[12][8] ), .A1(out_new[8]), .S(N3462), .Z(n1512)
         );
  CMX2X2 U4397 ( .A0(\memory[12][7] ), .A1(out_new[7]), .S(N3462), .Z(n1513)
         );
  CMX2X2 U4398 ( .A0(\memory[12][6] ), .A1(out_new[6]), .S(N3462), .Z(n1514)
         );
  CMX2X2 U4399 ( .A0(\memory[12][5] ), .A1(out_new[5]), .S(N3462), .Z(n1515)
         );
  CMX2X2 U4400 ( .A0(\memory[12][4] ), .A1(out_new[4]), .S(N3462), .Z(n1516)
         );
  CMX2X2 U4401 ( .A0(\memory[12][3] ), .A1(out_new[3]), .S(N3462), .Z(n1517)
         );
  CMX2X2 U4402 ( .A0(\memory[12][2] ), .A1(out_new[2]), .S(N3462), .Z(n1518)
         );
  CMX2X2 U4403 ( .A0(\memory[12][1] ), .A1(out_new[1]), .S(N3462), .Z(n1519)
         );
  CMX2X2 U4404 ( .A0(\memory[12][0] ), .A1(out_new[0]), .S(N3462), .Z(n1520)
         );
  CMX2X2 U4405 ( .A0(\memory[11][63] ), .A1(out_new[63]), .S(N3391), .Z(n1528)
         );
  CMX2X2 U4406 ( .A0(\memory[11][62] ), .A1(out_new[62]), .S(N3391), .Z(n1529)
         );
  CMX2X2 U4407 ( .A0(\memory[11][61] ), .A1(out_new[61]), .S(N3391), .Z(n1530)
         );
  CMX2X2 U4408 ( .A0(\memory[11][60] ), .A1(out_new[60]), .S(N3391), .Z(n1531)
         );
  CMX2X2 U4409 ( .A0(\memory[11][59] ), .A1(out_new[59]), .S(N3391), .Z(n1532)
         );
  CMX2X2 U4410 ( .A0(\memory[11][58] ), .A1(out_new[58]), .S(N3391), .Z(n1533)
         );
  CMX2X2 U4411 ( .A0(\memory[11][57] ), .A1(out_new[57]), .S(N3391), .Z(n1534)
         );
  CMX2X2 U4412 ( .A0(\memory[11][56] ), .A1(out_new[56]), .S(N3391), .Z(n1535)
         );
  CMX2X2 U4413 ( .A0(\memory[11][55] ), .A1(out_new[55]), .S(N3391), .Z(n1536)
         );
  CMX2X2 U4414 ( .A0(\memory[11][54] ), .A1(out_new[54]), .S(N3391), .Z(n1537)
         );
  CMX2X2 U4415 ( .A0(\memory[11][53] ), .A1(out_new[53]), .S(N3391), .Z(n1538)
         );
  CMX2X2 U4416 ( .A0(\memory[11][52] ), .A1(out_new[52]), .S(N3391), .Z(n1539)
         );
  CMX2X2 U4417 ( .A0(\memory[11][51] ), .A1(out_new[51]), .S(N3391), .Z(n1540)
         );
  CMX2X2 U4418 ( .A0(\memory[11][50] ), .A1(out_new[50]), .S(N3391), .Z(n1541)
         );
  CMX2X2 U4419 ( .A0(\memory[11][49] ), .A1(out_new[49]), .S(N3391), .Z(n1542)
         );
  CMX2X2 U4420 ( .A0(\memory[11][48] ), .A1(out_new[48]), .S(N3391), .Z(n1543)
         );
  CMX2X2 U4421 ( .A0(\memory[11][47] ), .A1(out_new[47]), .S(N3391), .Z(n1544)
         );
  CMX2X2 U4422 ( .A0(\memory[11][46] ), .A1(out_new[46]), .S(N3391), .Z(n1545)
         );
  CMX2X2 U4423 ( .A0(\memory[11][45] ), .A1(out_new[45]), .S(N3391), .Z(n1546)
         );
  CMX2X2 U4424 ( .A0(\memory[11][44] ), .A1(out_new[44]), .S(N3391), .Z(n1547)
         );
  CMX2X2 U4425 ( .A0(\memory[11][43] ), .A1(out_new[43]), .S(N3391), .Z(n1548)
         );
  CMX2X2 U4426 ( .A0(\memory[11][42] ), .A1(out_new[42]), .S(N3391), .Z(n1549)
         );
  CMX2X2 U4427 ( .A0(\memory[11][41] ), .A1(out_new[41]), .S(N3391), .Z(n1550)
         );
  CMX2X2 U4428 ( .A0(\memory[11][40] ), .A1(out_new[40]), .S(N3391), .Z(n1551)
         );
  CMX2X2 U4429 ( .A0(\memory[11][39] ), .A1(out_new[39]), .S(N3391), .Z(n1552)
         );
  CMX2X2 U4430 ( .A0(\memory[11][38] ), .A1(out_new[38]), .S(N3391), .Z(n1553)
         );
  CMX2X2 U4431 ( .A0(\memory[11][37] ), .A1(out_new[37]), .S(N3391), .Z(n1554)
         );
  CMX2X2 U4432 ( .A0(\memory[11][36] ), .A1(out_new[36]), .S(N3391), .Z(n1555)
         );
  CMX2X2 U4433 ( .A0(\memory[11][35] ), .A1(out_new[35]), .S(N3391), .Z(n1556)
         );
  CMX2X2 U4434 ( .A0(\memory[11][34] ), .A1(out_new[34]), .S(N3391), .Z(n1557)
         );
  CMX2X2 U4435 ( .A0(\memory[11][33] ), .A1(out_new[33]), .S(N3391), .Z(n1558)
         );
  CMX2X2 U4436 ( .A0(\memory[11][32] ), .A1(out_new[32]), .S(N3391), .Z(n1559)
         );
  CMX2X2 U4437 ( .A0(\memory[11][31] ), .A1(out_new[31]), .S(N3391), .Z(n1560)
         );
  CMX2X2 U4438 ( .A0(\memory[11][30] ), .A1(out_new[30]), .S(N3391), .Z(n1561)
         );
  CMX2X2 U4439 ( .A0(\memory[11][29] ), .A1(out_new[29]), .S(N3391), .Z(n1562)
         );
  CMX2X2 U4440 ( .A0(\memory[11][28] ), .A1(out_new[28]), .S(N3391), .Z(n1563)
         );
  CMX2X2 U4441 ( .A0(\memory[11][27] ), .A1(out_new[27]), .S(N3391), .Z(n1564)
         );
  CMX2X2 U4442 ( .A0(\memory[11][26] ), .A1(out_new[26]), .S(N3391), .Z(n1565)
         );
  CMX2X2 U4443 ( .A0(\memory[11][25] ), .A1(out_new[25]), .S(N3391), .Z(n1566)
         );
  CMX2X2 U4444 ( .A0(\memory[11][24] ), .A1(out_new[24]), .S(N3391), .Z(n1567)
         );
  CMX2X2 U4445 ( .A0(\memory[11][23] ), .A1(out_new[23]), .S(N3391), .Z(n1568)
         );
  CMX2X2 U4446 ( .A0(\memory[11][22] ), .A1(out_new[22]), .S(N3391), .Z(n1569)
         );
  CMX2X2 U4447 ( .A0(\memory[11][21] ), .A1(out_new[21]), .S(N3391), .Z(n1570)
         );
  CMX2X2 U4448 ( .A0(\memory[11][20] ), .A1(out_new[20]), .S(N3391), .Z(n1571)
         );
  CMX2X2 U4449 ( .A0(\memory[11][19] ), .A1(out_new[19]), .S(N3391), .Z(n1572)
         );
  CMX2X2 U4450 ( .A0(\memory[11][18] ), .A1(out_new[18]), .S(N3391), .Z(n1573)
         );
  CMX2X2 U4451 ( .A0(\memory[11][17] ), .A1(out_new[17]), .S(N3391), .Z(n1574)
         );
  CMX2X2 U4452 ( .A0(\memory[11][16] ), .A1(out_new[16]), .S(N3391), .Z(n1575)
         );
  CMX2X2 U4453 ( .A0(\memory[11][15] ), .A1(out_new[15]), .S(N3391), .Z(n1576)
         );
  CMX2X2 U4454 ( .A0(\memory[11][14] ), .A1(out_new[14]), .S(N3391), .Z(n1577)
         );
  CMX2X2 U4455 ( .A0(\memory[11][13] ), .A1(out_new[13]), .S(N3391), .Z(n1578)
         );
  CMX2X2 U4456 ( .A0(\memory[11][12] ), .A1(out_new[12]), .S(N3391), .Z(n1579)
         );
  CMX2X2 U4457 ( .A0(\memory[11][11] ), .A1(out_new[11]), .S(N3391), .Z(n1580)
         );
  CMX2X2 U4458 ( .A0(\memory[11][10] ), .A1(out_new[10]), .S(N3391), .Z(n1581)
         );
  CMX2X2 U4459 ( .A0(\memory[11][9] ), .A1(out_new[9]), .S(N3391), .Z(n1582)
         );
  CMX2X2 U4460 ( .A0(\memory[11][8] ), .A1(out_new[8]), .S(N3391), .Z(n1583)
         );
  CMX2X2 U4461 ( .A0(\memory[11][7] ), .A1(out_new[7]), .S(N3391), .Z(n1584)
         );
  CMX2X2 U4462 ( .A0(\memory[11][6] ), .A1(out_new[6]), .S(N3391), .Z(n1585)
         );
  CMX2X2 U4463 ( .A0(\memory[11][5] ), .A1(out_new[5]), .S(N3391), .Z(n1586)
         );
  CMX2X2 U4464 ( .A0(\memory[11][4] ), .A1(out_new[4]), .S(N3391), .Z(n1587)
         );
  CMX2X2 U4465 ( .A0(\memory[11][3] ), .A1(out_new[3]), .S(N3391), .Z(n1588)
         );
  CMX2X2 U4466 ( .A0(\memory[11][2] ), .A1(out_new[2]), .S(N3391), .Z(n1589)
         );
  CMX2X2 U4467 ( .A0(\memory[11][1] ), .A1(out_new[1]), .S(N3391), .Z(n1590)
         );
  CMX2X2 U4468 ( .A0(\memory[11][0] ), .A1(out_new[0]), .S(N3391), .Z(n1591)
         );
  CMX2X2 U4469 ( .A0(\memory[10][63] ), .A1(out_new[63]), .S(N3320), .Z(n1599)
         );
  CMX2X2 U4470 ( .A0(\memory[10][62] ), .A1(out_new[62]), .S(N3320), .Z(n1600)
         );
  CMX2X2 U4471 ( .A0(\memory[10][61] ), .A1(out_new[61]), .S(N3320), .Z(n1601)
         );
  CMX2X2 U4472 ( .A0(\memory[10][60] ), .A1(out_new[60]), .S(N3320), .Z(n1602)
         );
  CMX2X2 U4473 ( .A0(\memory[10][59] ), .A1(out_new[59]), .S(N3320), .Z(n1603)
         );
  CMX2X2 U4474 ( .A0(\memory[10][58] ), .A1(out_new[58]), .S(N3320), .Z(n1604)
         );
  CMX2X2 U4475 ( .A0(\memory[10][57] ), .A1(out_new[57]), .S(N3320), .Z(n1605)
         );
  CMX2X2 U4476 ( .A0(\memory[10][56] ), .A1(out_new[56]), .S(N3320), .Z(n1606)
         );
  CMX2X2 U4477 ( .A0(\memory[10][55] ), .A1(out_new[55]), .S(N3320), .Z(n1607)
         );
  CMX2X2 U4478 ( .A0(\memory[10][54] ), .A1(out_new[54]), .S(N3320), .Z(n1608)
         );
  CMX2X2 U4479 ( .A0(\memory[10][53] ), .A1(out_new[53]), .S(N3320), .Z(n1609)
         );
  CMX2X2 U4480 ( .A0(\memory[10][52] ), .A1(out_new[52]), .S(N3320), .Z(n1610)
         );
  CMX2X2 U4481 ( .A0(\memory[10][51] ), .A1(out_new[51]), .S(N3320), .Z(n1611)
         );
  CMX2X2 U4482 ( .A0(\memory[10][50] ), .A1(out_new[50]), .S(N3320), .Z(n1612)
         );
  CMX2X2 U4483 ( .A0(\memory[10][49] ), .A1(out_new[49]), .S(N3320), .Z(n1613)
         );
  CMX2X2 U4484 ( .A0(\memory[10][48] ), .A1(out_new[48]), .S(N3320), .Z(n1614)
         );
  CMX2X2 U4485 ( .A0(\memory[10][47] ), .A1(out_new[47]), .S(N3320), .Z(n1615)
         );
  CMX2X2 U4486 ( .A0(\memory[10][46] ), .A1(out_new[46]), .S(N3320), .Z(n1616)
         );
  CMX2X2 U4487 ( .A0(\memory[10][45] ), .A1(out_new[45]), .S(N3320), .Z(n1617)
         );
  CMX2X2 U4488 ( .A0(\memory[10][44] ), .A1(out_new[44]), .S(N3320), .Z(n1618)
         );
  CMX2X2 U4489 ( .A0(\memory[10][43] ), .A1(out_new[43]), .S(N3320), .Z(n1619)
         );
  CMX2X2 U4490 ( .A0(\memory[10][42] ), .A1(out_new[42]), .S(N3320), .Z(n1620)
         );
  CMX2X2 U4491 ( .A0(\memory[10][41] ), .A1(out_new[41]), .S(N3320), .Z(n1621)
         );
  CMX2X2 U4492 ( .A0(\memory[10][40] ), .A1(out_new[40]), .S(N3320), .Z(n1622)
         );
  CMX2X2 U4493 ( .A0(\memory[10][39] ), .A1(out_new[39]), .S(N3320), .Z(n1623)
         );
  CMX2X2 U4494 ( .A0(\memory[10][38] ), .A1(out_new[38]), .S(N3320), .Z(n1624)
         );
  CMX2X2 U4495 ( .A0(\memory[10][37] ), .A1(out_new[37]), .S(N3320), .Z(n1625)
         );
  CMX2X2 U4496 ( .A0(\memory[10][36] ), .A1(out_new[36]), .S(N3320), .Z(n1626)
         );
  CMX2X2 U4497 ( .A0(\memory[10][35] ), .A1(out_new[35]), .S(N3320), .Z(n1627)
         );
  CMX2X2 U4498 ( .A0(\memory[10][34] ), .A1(out_new[34]), .S(N3320), .Z(n1628)
         );
  CMX2X2 U4499 ( .A0(\memory[10][33] ), .A1(out_new[33]), .S(N3320), .Z(n1629)
         );
  CMX2X2 U4500 ( .A0(\memory[10][32] ), .A1(out_new[32]), .S(N3320), .Z(n1630)
         );
  CMX2X2 U4501 ( .A0(\memory[10][31] ), .A1(out_new[31]), .S(N3320), .Z(n1631)
         );
  CMX2X2 U4502 ( .A0(\memory[10][30] ), .A1(out_new[30]), .S(N3320), .Z(n1632)
         );
  CMX2X2 U4503 ( .A0(\memory[10][29] ), .A1(out_new[29]), .S(N3320), .Z(n1633)
         );
  CMX2X2 U4504 ( .A0(\memory[10][28] ), .A1(out_new[28]), .S(N3320), .Z(n1634)
         );
  CMX2X2 U4505 ( .A0(\memory[10][27] ), .A1(out_new[27]), .S(N3320), .Z(n1635)
         );
  CMX2X2 U4506 ( .A0(\memory[10][26] ), .A1(out_new[26]), .S(N3320), .Z(n1636)
         );
  CMX2X2 U4507 ( .A0(\memory[10][25] ), .A1(out_new[25]), .S(N3320), .Z(n1637)
         );
  CMX2X2 U4508 ( .A0(\memory[10][24] ), .A1(out_new[24]), .S(N3320), .Z(n1638)
         );
  CMX2X2 U4509 ( .A0(\memory[10][23] ), .A1(out_new[23]), .S(N3320), .Z(n1639)
         );
  CMX2X2 U4510 ( .A0(\memory[10][22] ), .A1(out_new[22]), .S(N3320), .Z(n1640)
         );
  CMX2X2 U4511 ( .A0(\memory[10][21] ), .A1(out_new[21]), .S(N3320), .Z(n1641)
         );
  CMX2X2 U4512 ( .A0(\memory[10][20] ), .A1(out_new[20]), .S(N3320), .Z(n1642)
         );
  CMX2X2 U4513 ( .A0(\memory[10][19] ), .A1(out_new[19]), .S(N3320), .Z(n1643)
         );
  CMX2X2 U4514 ( .A0(\memory[10][18] ), .A1(out_new[18]), .S(N3320), .Z(n1644)
         );
  CMX2X2 U4515 ( .A0(\memory[10][17] ), .A1(out_new[17]), .S(N3320), .Z(n1645)
         );
  CMX2X2 U4516 ( .A0(\memory[10][16] ), .A1(out_new[16]), .S(N3320), .Z(n1646)
         );
  CMX2X2 U4517 ( .A0(\memory[10][15] ), .A1(out_new[15]), .S(N3320), .Z(n1647)
         );
  CMX2X2 U4518 ( .A0(\memory[10][14] ), .A1(out_new[14]), .S(N3320), .Z(n1648)
         );
  CMX2X2 U4519 ( .A0(\memory[10][13] ), .A1(out_new[13]), .S(N3320), .Z(n1649)
         );
  CMX2X2 U4520 ( .A0(\memory[10][12] ), .A1(out_new[12]), .S(N3320), .Z(n1650)
         );
  CMX2X2 U4521 ( .A0(\memory[10][11] ), .A1(out_new[11]), .S(N3320), .Z(n1651)
         );
  CMX2X2 U4522 ( .A0(\memory[10][10] ), .A1(out_new[10]), .S(N3320), .Z(n1652)
         );
  CMX2X2 U4523 ( .A0(\memory[10][9] ), .A1(out_new[9]), .S(N3320), .Z(n1653)
         );
  CMX2X2 U4524 ( .A0(\memory[10][8] ), .A1(out_new[8]), .S(N3320), .Z(n1654)
         );
  CMX2X2 U4525 ( .A0(\memory[10][7] ), .A1(out_new[7]), .S(N3320), .Z(n1655)
         );
  CMX2X2 U4526 ( .A0(\memory[10][6] ), .A1(out_new[6]), .S(N3320), .Z(n1656)
         );
  CMX2X2 U4527 ( .A0(\memory[10][5] ), .A1(out_new[5]), .S(N3320), .Z(n1657)
         );
  CMX2X2 U4528 ( .A0(\memory[10][4] ), .A1(out_new[4]), .S(N3320), .Z(n1658)
         );
  CMX2X2 U4529 ( .A0(\memory[10][3] ), .A1(out_new[3]), .S(N3320), .Z(n1659)
         );
  CMX2X2 U4530 ( .A0(\memory[10][2] ), .A1(out_new[2]), .S(N3320), .Z(n1660)
         );
  CMX2X2 U4531 ( .A0(\memory[10][1] ), .A1(out_new[1]), .S(N3320), .Z(n1661)
         );
  CMX2X2 U4532 ( .A0(\memory[10][0] ), .A1(out_new[0]), .S(N3320), .Z(n1662)
         );
  CMX2X2 U4533 ( .A0(\memory[9][63] ), .A1(out_new[63]), .S(N3249), .Z(n1670)
         );
  CMX2X2 U4534 ( .A0(\memory[9][62] ), .A1(out_new[62]), .S(N3249), .Z(n1671)
         );
  CMX2X2 U4535 ( .A0(\memory[9][61] ), .A1(out_new[61]), .S(N3249), .Z(n1672)
         );
  CMX2X2 U4536 ( .A0(\memory[9][60] ), .A1(out_new[60]), .S(N3249), .Z(n1673)
         );
  CMX2X2 U4537 ( .A0(\memory[9][59] ), .A1(out_new[59]), .S(N3249), .Z(n1674)
         );
  CMX2X2 U4538 ( .A0(\memory[9][58] ), .A1(out_new[58]), .S(N3249), .Z(n1675)
         );
  CMX2X2 U4539 ( .A0(\memory[9][57] ), .A1(out_new[57]), .S(N3249), .Z(n1676)
         );
  CMX2X2 U4540 ( .A0(\memory[9][56] ), .A1(out_new[56]), .S(N3249), .Z(n1677)
         );
  CMX2X2 U4541 ( .A0(\memory[9][55] ), .A1(out_new[55]), .S(N3249), .Z(n1678)
         );
  CMX2X2 U4542 ( .A0(\memory[9][54] ), .A1(out_new[54]), .S(N3249), .Z(n1679)
         );
  CMX2X2 U4543 ( .A0(\memory[9][53] ), .A1(out_new[53]), .S(N3249), .Z(n1680)
         );
  CMX2X2 U4544 ( .A0(\memory[9][52] ), .A1(out_new[52]), .S(N3249), .Z(n1681)
         );
  CMX2X2 U4545 ( .A0(\memory[9][51] ), .A1(out_new[51]), .S(N3249), .Z(n1682)
         );
  CMX2X2 U4546 ( .A0(\memory[9][50] ), .A1(out_new[50]), .S(N3249), .Z(n1683)
         );
  CMX2X2 U4547 ( .A0(\memory[9][49] ), .A1(out_new[49]), .S(N3249), .Z(n1684)
         );
  CMX2X2 U4548 ( .A0(\memory[9][48] ), .A1(out_new[48]), .S(N3249), .Z(n1685)
         );
  CMX2X2 U4549 ( .A0(\memory[9][47] ), .A1(out_new[47]), .S(N3249), .Z(n1686)
         );
  CMX2X2 U4550 ( .A0(\memory[9][46] ), .A1(out_new[46]), .S(N3249), .Z(n1687)
         );
  CMX2X2 U4551 ( .A0(\memory[9][45] ), .A1(out_new[45]), .S(N3249), .Z(n1688)
         );
  CMX2X2 U4552 ( .A0(\memory[9][44] ), .A1(out_new[44]), .S(N3249), .Z(n1689)
         );
  CMX2X2 U4553 ( .A0(\memory[9][43] ), .A1(out_new[43]), .S(N3249), .Z(n1690)
         );
  CMX2X2 U4554 ( .A0(\memory[9][42] ), .A1(out_new[42]), .S(N3249), .Z(n1691)
         );
  CMX2X2 U4555 ( .A0(\memory[9][41] ), .A1(out_new[41]), .S(N3249), .Z(n1692)
         );
  CMX2X2 U4556 ( .A0(\memory[9][40] ), .A1(out_new[40]), .S(N3249), .Z(n1693)
         );
  CMX2X2 U4557 ( .A0(\memory[9][39] ), .A1(out_new[39]), .S(N3249), .Z(n1694)
         );
  CMX2X2 U4558 ( .A0(\memory[9][38] ), .A1(out_new[38]), .S(N3249), .Z(n1695)
         );
  CMX2X2 U4559 ( .A0(\memory[9][37] ), .A1(out_new[37]), .S(N3249), .Z(n1696)
         );
  CMX2X2 U4560 ( .A0(\memory[9][36] ), .A1(out_new[36]), .S(N3249), .Z(n1697)
         );
  CMX2X2 U4561 ( .A0(\memory[9][35] ), .A1(out_new[35]), .S(N3249), .Z(n1698)
         );
  CMX2X2 U4562 ( .A0(\memory[9][34] ), .A1(out_new[34]), .S(N3249), .Z(n1699)
         );
  CMX2X2 U4563 ( .A0(\memory[9][33] ), .A1(out_new[33]), .S(N3249), .Z(n1700)
         );
  CMX2X2 U4564 ( .A0(\memory[9][32] ), .A1(out_new[32]), .S(N3249), .Z(n1701)
         );
  CMX2X2 U4565 ( .A0(\memory[9][31] ), .A1(out_new[31]), .S(N3249), .Z(n1702)
         );
  CMX2X2 U4566 ( .A0(\memory[9][30] ), .A1(out_new[30]), .S(N3249), .Z(n1703)
         );
  CMX2X2 U4567 ( .A0(\memory[9][29] ), .A1(out_new[29]), .S(N3249), .Z(n1704)
         );
  CMX2X2 U4568 ( .A0(\memory[9][28] ), .A1(out_new[28]), .S(N3249), .Z(n1705)
         );
  CMX2X2 U4569 ( .A0(\memory[9][27] ), .A1(out_new[27]), .S(N3249), .Z(n1706)
         );
  CMX2X2 U4570 ( .A0(\memory[9][26] ), .A1(out_new[26]), .S(N3249), .Z(n1707)
         );
  CMX2X2 U4571 ( .A0(\memory[9][25] ), .A1(out_new[25]), .S(N3249), .Z(n1708)
         );
  CMX2X2 U4572 ( .A0(\memory[9][24] ), .A1(out_new[24]), .S(N3249), .Z(n1709)
         );
  CMX2X2 U4573 ( .A0(\memory[9][23] ), .A1(out_new[23]), .S(N3249), .Z(n1710)
         );
  CMX2X2 U4574 ( .A0(\memory[9][22] ), .A1(out_new[22]), .S(N3249), .Z(n1711)
         );
  CMX2X2 U4575 ( .A0(\memory[9][21] ), .A1(out_new[21]), .S(N3249), .Z(n1712)
         );
  CMX2X2 U4576 ( .A0(\memory[9][20] ), .A1(out_new[20]), .S(N3249), .Z(n1713)
         );
  CMX2X2 U4577 ( .A0(\memory[9][19] ), .A1(out_new[19]), .S(N3249), .Z(n1714)
         );
  CMX2X2 U4578 ( .A0(\memory[9][18] ), .A1(out_new[18]), .S(N3249), .Z(n1715)
         );
  CMX2X2 U4579 ( .A0(\memory[9][17] ), .A1(out_new[17]), .S(N3249), .Z(n1716)
         );
  CMX2X2 U4580 ( .A0(\memory[9][16] ), .A1(out_new[16]), .S(N3249), .Z(n1717)
         );
  CMX2X2 U4581 ( .A0(\memory[9][15] ), .A1(out_new[15]), .S(N3249), .Z(n1718)
         );
  CMX2X2 U4582 ( .A0(\memory[9][14] ), .A1(out_new[14]), .S(N3249), .Z(n1719)
         );
  CMX2X2 U4583 ( .A0(\memory[9][13] ), .A1(out_new[13]), .S(N3249), .Z(n1720)
         );
  CMX2X2 U4584 ( .A0(\memory[9][12] ), .A1(out_new[12]), .S(N3249), .Z(n1721)
         );
  CMX2X2 U4585 ( .A0(\memory[9][11] ), .A1(out_new[11]), .S(N3249), .Z(n1722)
         );
  CMX2X2 U4586 ( .A0(\memory[9][10] ), .A1(out_new[10]), .S(N3249), .Z(n1723)
         );
  CMX2X2 U4587 ( .A0(\memory[9][9] ), .A1(out_new[9]), .S(N3249), .Z(n1724) );
  CMX2X2 U4588 ( .A0(\memory[9][8] ), .A1(out_new[8]), .S(N3249), .Z(n1725) );
  CMX2X2 U4589 ( .A0(\memory[9][7] ), .A1(out_new[7]), .S(N3249), .Z(n1726) );
  CMX2X2 U4590 ( .A0(\memory[9][6] ), .A1(out_new[6]), .S(N3249), .Z(n1727) );
  CMX2X2 U4591 ( .A0(\memory[9][5] ), .A1(out_new[5]), .S(N3249), .Z(n1728) );
  CMX2X2 U4592 ( .A0(\memory[9][4] ), .A1(out_new[4]), .S(N3249), .Z(n1729) );
  CMX2X2 U4593 ( .A0(\memory[9][3] ), .A1(out_new[3]), .S(N3249), .Z(n1730) );
  CMX2X2 U4594 ( .A0(\memory[9][2] ), .A1(out_new[2]), .S(N3249), .Z(n1731) );
  CMX2X2 U4595 ( .A0(\memory[9][1] ), .A1(out_new[1]), .S(N3249), .Z(n1732) );
  CMX2X2 U4596 ( .A0(\memory[9][0] ), .A1(out_new[0]), .S(N3249), .Z(n1733) );
  CMX2X2 U4597 ( .A0(\memory[8][63] ), .A1(out_new[63]), .S(N3178), .Z(n1741)
         );
  CMX2X2 U4598 ( .A0(\memory[8][62] ), .A1(out_new[62]), .S(N3178), .Z(n1742)
         );
  CMX2X2 U4599 ( .A0(\memory[8][61] ), .A1(out_new[61]), .S(N3178), .Z(n1743)
         );
  CMX2X2 U4600 ( .A0(\memory[8][60] ), .A1(out_new[60]), .S(N3178), .Z(n1744)
         );
  CMX2X2 U4601 ( .A0(\memory[8][59] ), .A1(out_new[59]), .S(N3178), .Z(n1745)
         );
  CMX2X2 U4602 ( .A0(\memory[8][58] ), .A1(out_new[58]), .S(N3178), .Z(n1746)
         );
  CMX2X2 U4603 ( .A0(\memory[8][57] ), .A1(out_new[57]), .S(N3178), .Z(n1747)
         );
  CMX2X2 U4604 ( .A0(\memory[8][56] ), .A1(out_new[56]), .S(N3178), .Z(n1748)
         );
  CMX2X2 U4605 ( .A0(\memory[8][55] ), .A1(out_new[55]), .S(N3178), .Z(n1749)
         );
  CMX2X2 U4606 ( .A0(\memory[8][54] ), .A1(out_new[54]), .S(N3178), .Z(n1750)
         );
  CMX2X2 U4607 ( .A0(\memory[8][53] ), .A1(out_new[53]), .S(N3178), .Z(n1751)
         );
  CMX2X2 U4608 ( .A0(\memory[8][52] ), .A1(out_new[52]), .S(N3178), .Z(n1752)
         );
  CMX2X2 U4609 ( .A0(\memory[8][51] ), .A1(out_new[51]), .S(N3178), .Z(n1753)
         );
  CMX2X2 U4610 ( .A0(\memory[8][50] ), .A1(out_new[50]), .S(N3178), .Z(n1754)
         );
  CMX2X2 U4611 ( .A0(\memory[8][49] ), .A1(out_new[49]), .S(N3178), .Z(n1755)
         );
  CMX2X2 U4612 ( .A0(\memory[8][48] ), .A1(out_new[48]), .S(N3178), .Z(n1756)
         );
  CMX2X2 U4613 ( .A0(\memory[8][47] ), .A1(out_new[47]), .S(N3178), .Z(n1757)
         );
  CMX2X2 U4614 ( .A0(\memory[8][46] ), .A1(out_new[46]), .S(N3178), .Z(n1758)
         );
  CMX2X2 U4615 ( .A0(\memory[8][45] ), .A1(out_new[45]), .S(N3178), .Z(n1759)
         );
  CMX2X2 U4616 ( .A0(\memory[8][44] ), .A1(out_new[44]), .S(N3178), .Z(n1760)
         );
  CMX2X2 U4617 ( .A0(\memory[8][43] ), .A1(out_new[43]), .S(N3178), .Z(n1761)
         );
  CMX2X2 U4618 ( .A0(\memory[8][42] ), .A1(out_new[42]), .S(N3178), .Z(n1762)
         );
  CMX2X2 U4619 ( .A0(\memory[8][41] ), .A1(out_new[41]), .S(N3178), .Z(n1763)
         );
  CMX2X2 U4620 ( .A0(\memory[8][40] ), .A1(out_new[40]), .S(N3178), .Z(n1764)
         );
  CMX2X2 U4621 ( .A0(\memory[8][39] ), .A1(out_new[39]), .S(N3178), .Z(n1765)
         );
  CMX2X2 U4622 ( .A0(\memory[8][38] ), .A1(out_new[38]), .S(N3178), .Z(n1766)
         );
  CMX2X2 U4623 ( .A0(\memory[8][37] ), .A1(out_new[37]), .S(N3178), .Z(n1767)
         );
  CMX2X2 U4624 ( .A0(\memory[8][36] ), .A1(out_new[36]), .S(N3178), .Z(n1768)
         );
  CMX2X2 U4625 ( .A0(\memory[8][35] ), .A1(out_new[35]), .S(N3178), .Z(n1769)
         );
  CMX2X2 U4626 ( .A0(\memory[8][34] ), .A1(out_new[34]), .S(N3178), .Z(n1770)
         );
  CMX2X2 U4627 ( .A0(\memory[8][33] ), .A1(out_new[33]), .S(N3178), .Z(n1771)
         );
  CMX2X2 U4628 ( .A0(\memory[8][32] ), .A1(out_new[32]), .S(N3178), .Z(n1772)
         );
  CMX2X2 U4629 ( .A0(\memory[8][31] ), .A1(out_new[31]), .S(N3178), .Z(n1773)
         );
  CMX2X2 U4630 ( .A0(\memory[8][30] ), .A1(out_new[30]), .S(N3178), .Z(n1774)
         );
  CMX2X2 U4631 ( .A0(\memory[8][29] ), .A1(out_new[29]), .S(N3178), .Z(n1775)
         );
  CMX2X2 U4632 ( .A0(\memory[8][28] ), .A1(out_new[28]), .S(N3178), .Z(n1776)
         );
  CMX2X2 U4633 ( .A0(\memory[8][27] ), .A1(out_new[27]), .S(N3178), .Z(n1777)
         );
  CMX2X2 U4634 ( .A0(\memory[8][26] ), .A1(out_new[26]), .S(N3178), .Z(n1778)
         );
  CMX2X2 U4635 ( .A0(\memory[8][25] ), .A1(out_new[25]), .S(N3178), .Z(n1779)
         );
  CMX2X2 U4636 ( .A0(\memory[8][24] ), .A1(out_new[24]), .S(N3178), .Z(n1780)
         );
  CMX2X2 U4637 ( .A0(\memory[8][23] ), .A1(out_new[23]), .S(N3178), .Z(n1781)
         );
  CMX2X2 U4638 ( .A0(\memory[8][22] ), .A1(out_new[22]), .S(N3178), .Z(n1782)
         );
  CMX2X2 U4639 ( .A0(\memory[8][21] ), .A1(out_new[21]), .S(N3178), .Z(n1783)
         );
  CMX2X2 U4640 ( .A0(\memory[8][20] ), .A1(out_new[20]), .S(N3178), .Z(n1784)
         );
  CMX2X2 U4641 ( .A0(\memory[8][19] ), .A1(out_new[19]), .S(N3178), .Z(n1785)
         );
  CMX2X2 U4642 ( .A0(\memory[8][18] ), .A1(out_new[18]), .S(N3178), .Z(n1786)
         );
  CMX2X2 U4643 ( .A0(\memory[8][17] ), .A1(out_new[17]), .S(N3178), .Z(n1787)
         );
  CMX2X2 U4644 ( .A0(\memory[8][16] ), .A1(out_new[16]), .S(N3178), .Z(n1788)
         );
  CMX2X2 U4645 ( .A0(\memory[8][15] ), .A1(out_new[15]), .S(N3178), .Z(n1789)
         );
  CMX2X2 U4646 ( .A0(\memory[8][14] ), .A1(out_new[14]), .S(N3178), .Z(n1790)
         );
  CMX2X2 U4647 ( .A0(\memory[8][13] ), .A1(out_new[13]), .S(N3178), .Z(n1791)
         );
  CMX2X2 U4648 ( .A0(\memory[8][12] ), .A1(out_new[12]), .S(N3178), .Z(n1792)
         );
  CMX2X2 U4649 ( .A0(\memory[8][11] ), .A1(out_new[11]), .S(N3178), .Z(n1793)
         );
  CMX2X2 U4650 ( .A0(\memory[8][10] ), .A1(out_new[10]), .S(N3178), .Z(n1794)
         );
  CMX2X2 U4651 ( .A0(\memory[8][9] ), .A1(out_new[9]), .S(N3178), .Z(n1795) );
  CMX2X2 U4652 ( .A0(\memory[8][8] ), .A1(out_new[8]), .S(N3178), .Z(n1796) );
  CMX2X2 U4653 ( .A0(\memory[8][7] ), .A1(out_new[7]), .S(N3178), .Z(n1797) );
  CMX2X2 U4654 ( .A0(\memory[8][6] ), .A1(out_new[6]), .S(N3178), .Z(n1798) );
  CMX2X2 U4655 ( .A0(\memory[8][5] ), .A1(out_new[5]), .S(N3178), .Z(n1799) );
  CMX2X2 U4656 ( .A0(\memory[8][4] ), .A1(out_new[4]), .S(N3178), .Z(n1800) );
  CMX2X2 U4657 ( .A0(\memory[8][3] ), .A1(out_new[3]), .S(N3178), .Z(n1801) );
  CMX2X2 U4658 ( .A0(\memory[8][2] ), .A1(out_new[2]), .S(N3178), .Z(n1802) );
  CMX2X2 U4659 ( .A0(\memory[8][1] ), .A1(out_new[1]), .S(N3178), .Z(n1803) );
  CMX2X2 U4660 ( .A0(\memory[8][0] ), .A1(out_new[0]), .S(N3178), .Z(n1804) );
  CMX2X2 U4661 ( .A0(\memory[6][63] ), .A1(out_new[63]), .S(N3036), .Z(n1883)
         );
  CMX2X2 U4662 ( .A0(\memory[6][62] ), .A1(out_new[62]), .S(N3036), .Z(n1884)
         );
  CMX2X2 U4663 ( .A0(\memory[6][61] ), .A1(out_new[61]), .S(N3036), .Z(n1885)
         );
  CMX2X2 U4664 ( .A0(\memory[6][60] ), .A1(out_new[60]), .S(N3036), .Z(n1886)
         );
  CMX2X2 U4665 ( .A0(\memory[6][59] ), .A1(out_new[59]), .S(N3036), .Z(n1887)
         );
  CMX2X2 U4666 ( .A0(\memory[6][58] ), .A1(out_new[58]), .S(N3036), .Z(n1888)
         );
  CMX2X2 U4667 ( .A0(\memory[6][57] ), .A1(out_new[57]), .S(N3036), .Z(n1889)
         );
  CMX2X2 U4668 ( .A0(\memory[6][56] ), .A1(out_new[56]), .S(N3036), .Z(n1890)
         );
  CMX2X2 U4669 ( .A0(\memory[6][55] ), .A1(out_new[55]), .S(N3036), .Z(n1891)
         );
  CMX2X2 U4670 ( .A0(\memory[6][54] ), .A1(out_new[54]), .S(N3036), .Z(n1892)
         );
  CMX2X2 U4671 ( .A0(\memory[6][53] ), .A1(out_new[53]), .S(N3036), .Z(n1893)
         );
  CMX2X2 U4672 ( .A0(\memory[6][52] ), .A1(out_new[52]), .S(N3036), .Z(n1894)
         );
  CMX2X2 U4673 ( .A0(\memory[6][51] ), .A1(out_new[51]), .S(N3036), .Z(n1895)
         );
  CMX2X2 U4674 ( .A0(\memory[6][50] ), .A1(out_new[50]), .S(N3036), .Z(n1896)
         );
  CMX2X2 U4675 ( .A0(\memory[6][49] ), .A1(out_new[49]), .S(N3036), .Z(n1897)
         );
  CMX2X2 U4676 ( .A0(\memory[6][48] ), .A1(out_new[48]), .S(N3036), .Z(n1898)
         );
  CMX2X2 U4677 ( .A0(\memory[6][47] ), .A1(out_new[47]), .S(N3036), .Z(n1899)
         );
  CMX2X2 U4678 ( .A0(\memory[6][46] ), .A1(out_new[46]), .S(N3036), .Z(n1900)
         );
  CMX2X2 U4679 ( .A0(\memory[6][45] ), .A1(out_new[45]), .S(N3036), .Z(n1901)
         );
  CMX2X2 U4680 ( .A0(\memory[6][44] ), .A1(out_new[44]), .S(N3036), .Z(n1902)
         );
  CMX2X2 U4681 ( .A0(\memory[6][43] ), .A1(out_new[43]), .S(N3036), .Z(n1903)
         );
  CMX2X2 U4682 ( .A0(\memory[6][42] ), .A1(out_new[42]), .S(N3036), .Z(n1904)
         );
  CMX2X2 U4683 ( .A0(\memory[6][41] ), .A1(out_new[41]), .S(N3036), .Z(n1905)
         );
  CMX2X2 U4684 ( .A0(\memory[6][40] ), .A1(out_new[40]), .S(N3036), .Z(n1906)
         );
  CMX2X2 U4685 ( .A0(\memory[6][39] ), .A1(out_new[39]), .S(N3036), .Z(n1907)
         );
  CMX2X2 U4686 ( .A0(\memory[6][38] ), .A1(out_new[38]), .S(N3036), .Z(n1908)
         );
  CMX2X2 U4687 ( .A0(\memory[6][37] ), .A1(out_new[37]), .S(N3036), .Z(n1909)
         );
  CMX2X2 U4688 ( .A0(\memory[6][36] ), .A1(out_new[36]), .S(N3036), .Z(n1910)
         );
  CMX2X2 U4689 ( .A0(\memory[6][35] ), .A1(out_new[35]), .S(N3036), .Z(n1911)
         );
  CMX2X2 U4690 ( .A0(\memory[6][34] ), .A1(out_new[34]), .S(N3036), .Z(n1912)
         );
  CMX2X2 U4691 ( .A0(\memory[6][33] ), .A1(out_new[33]), .S(N3036), .Z(n1913)
         );
  CMX2X2 U4692 ( .A0(\memory[6][32] ), .A1(out_new[32]), .S(N3036), .Z(n1914)
         );
  CMX2X2 U4693 ( .A0(\memory[6][31] ), .A1(out_new[31]), .S(N3036), .Z(n1915)
         );
  CMX2X2 U4694 ( .A0(\memory[6][30] ), .A1(out_new[30]), .S(N3036), .Z(n1916)
         );
  CMX2X2 U4695 ( .A0(\memory[6][29] ), .A1(out_new[29]), .S(N3036), .Z(n1917)
         );
  CMX2X2 U4696 ( .A0(\memory[6][28] ), .A1(out_new[28]), .S(N3036), .Z(n1918)
         );
  CMX2X2 U4697 ( .A0(\memory[6][27] ), .A1(out_new[27]), .S(N3036), .Z(n1919)
         );
  CMX2X2 U4698 ( .A0(\memory[6][26] ), .A1(out_new[26]), .S(N3036), .Z(n1920)
         );
  CMX2X2 U4699 ( .A0(\memory[6][25] ), .A1(out_new[25]), .S(N3036), .Z(n1921)
         );
  CMX2X2 U4700 ( .A0(\memory[6][24] ), .A1(out_new[24]), .S(N3036), .Z(n1922)
         );
  CMX2X2 U4701 ( .A0(\memory[6][23] ), .A1(out_new[23]), .S(N3036), .Z(n1923)
         );
  CMX2X2 U4702 ( .A0(\memory[6][22] ), .A1(out_new[22]), .S(N3036), .Z(n1924)
         );
  CMX2X2 U4703 ( .A0(\memory[6][21] ), .A1(out_new[21]), .S(N3036), .Z(n1925)
         );
  CMX2X2 U4704 ( .A0(\memory[6][20] ), .A1(out_new[20]), .S(N3036), .Z(n1926)
         );
  CMX2X2 U4705 ( .A0(\memory[6][19] ), .A1(out_new[19]), .S(N3036), .Z(n1927)
         );
  CMX2X2 U4706 ( .A0(\memory[6][18] ), .A1(out_new[18]), .S(N3036), .Z(n1928)
         );
  CMX2X2 U4707 ( .A0(\memory[6][17] ), .A1(out_new[17]), .S(N3036), .Z(n1929)
         );
  CMX2X2 U4708 ( .A0(\memory[6][16] ), .A1(out_new[16]), .S(N3036), .Z(n1930)
         );
  CMX2X2 U4709 ( .A0(\memory[6][15] ), .A1(out_new[15]), .S(N3036), .Z(n1931)
         );
  CMX2X2 U4710 ( .A0(\memory[6][14] ), .A1(out_new[14]), .S(N3036), .Z(n1932)
         );
  CMX2X2 U4711 ( .A0(\memory[6][13] ), .A1(out_new[13]), .S(N3036), .Z(n1933)
         );
  CMX2X2 U4712 ( .A0(\memory[6][12] ), .A1(out_new[12]), .S(N3036), .Z(n1934)
         );
  CMX2X2 U4713 ( .A0(\memory[6][11] ), .A1(out_new[11]), .S(N3036), .Z(n1935)
         );
  CMX2X2 U4714 ( .A0(\memory[6][10] ), .A1(out_new[10]), .S(N3036), .Z(n1936)
         );
  CMX2X2 U4715 ( .A0(\memory[6][9] ), .A1(out_new[9]), .S(N3036), .Z(n1937) );
  CMX2X2 U4716 ( .A0(\memory[6][8] ), .A1(out_new[8]), .S(N3036), .Z(n1938) );
  CMX2X2 U4717 ( .A0(\memory[6][7] ), .A1(out_new[7]), .S(N3036), .Z(n1939) );
  CMX2X2 U4718 ( .A0(\memory[6][6] ), .A1(out_new[6]), .S(N3036), .Z(n1940) );
  CMX2X2 U4719 ( .A0(\memory[6][5] ), .A1(out_new[5]), .S(N3036), .Z(n1941) );
  CMX2X2 U4720 ( .A0(\memory[6][4] ), .A1(out_new[4]), .S(N3036), .Z(n1942) );
  CMX2X2 U4721 ( .A0(\memory[6][3] ), .A1(out_new[3]), .S(N3036), .Z(n1943) );
  CMX2X2 U4722 ( .A0(\memory[6][2] ), .A1(out_new[2]), .S(N3036), .Z(n1944) );
  CMX2X2 U4723 ( .A0(\memory[6][1] ), .A1(out_new[1]), .S(N3036), .Z(n1945) );
  CMX2X2 U4724 ( .A0(\memory[6][0] ), .A1(out_new[0]), .S(N3036), .Z(n1946) );
  CMX2X4 U4725 ( .A0(\memory[5][63] ), .A1(out_new[63]), .S(N2965), .Z(n1954)
         );
  CMX2X4 U4726 ( .A0(\memory[5][62] ), .A1(out_new[62]), .S(N2965), .Z(n1955)
         );
  CMX2X4 U4727 ( .A0(\memory[5][61] ), .A1(out_new[61]), .S(N2965), .Z(n1956)
         );
  CMX2X4 U4728 ( .A0(\memory[5][60] ), .A1(out_new[60]), .S(N2965), .Z(n1957)
         );
  CMX2X4 U4729 ( .A0(\memory[5][59] ), .A1(out_new[59]), .S(N2965), .Z(n1958)
         );
  CMX2X4 U4730 ( .A0(\memory[5][58] ), .A1(out_new[58]), .S(N2965), .Z(n1959)
         );
  CMX2X4 U4731 ( .A0(\memory[5][57] ), .A1(out_new[57]), .S(N2965), .Z(n1960)
         );
  CMX2X4 U4732 ( .A0(\memory[5][56] ), .A1(out_new[56]), .S(N2965), .Z(n1961)
         );
  CMX2X4 U4733 ( .A0(\memory[5][55] ), .A1(out_new[55]), .S(N2965), .Z(n1962)
         );
  CMX2X4 U4734 ( .A0(\memory[5][54] ), .A1(out_new[54]), .S(N2965), .Z(n1963)
         );
  CMX2X4 U4735 ( .A0(\memory[5][53] ), .A1(out_new[53]), .S(N2965), .Z(n1964)
         );
  CMX2X4 U4736 ( .A0(\memory[5][52] ), .A1(out_new[52]), .S(N2965), .Z(n1965)
         );
  CMX2X4 U4737 ( .A0(\memory[5][51] ), .A1(out_new[51]), .S(N2965), .Z(n1966)
         );
  CMX2X4 U4738 ( .A0(\memory[5][50] ), .A1(out_new[50]), .S(N2965), .Z(n1967)
         );
  CMX2X4 U4739 ( .A0(\memory[5][49] ), .A1(out_new[49]), .S(N2965), .Z(n1968)
         );
  CMX2X4 U4740 ( .A0(\memory[5][48] ), .A1(out_new[48]), .S(N2965), .Z(n1969)
         );
  CMX2X4 U4741 ( .A0(\memory[5][47] ), .A1(out_new[47]), .S(N2965), .Z(n1970)
         );
  CMX2X4 U4742 ( .A0(\memory[5][46] ), .A1(out_new[46]), .S(N2965), .Z(n1971)
         );
  CMX2X4 U4743 ( .A0(\memory[5][45] ), .A1(out_new[45]), .S(N2965), .Z(n1972)
         );
  CMX2X4 U4744 ( .A0(\memory[5][44] ), .A1(out_new[44]), .S(N2965), .Z(n1973)
         );
  CMX2X4 U4745 ( .A0(\memory[5][43] ), .A1(out_new[43]), .S(N2965), .Z(n1974)
         );
  CMX2X4 U4746 ( .A0(\memory[5][42] ), .A1(out_new[42]), .S(N2965), .Z(n1975)
         );
  CMX2X4 U4747 ( .A0(\memory[5][41] ), .A1(out_new[41]), .S(N2965), .Z(n1976)
         );
  CMX2X4 U4748 ( .A0(\memory[5][40] ), .A1(out_new[40]), .S(N2965), .Z(n1977)
         );
  CMX2X4 U4749 ( .A0(\memory[5][39] ), .A1(out_new[39]), .S(N2965), .Z(n1978)
         );
  CMX2X4 U4750 ( .A0(\memory[5][38] ), .A1(out_new[38]), .S(N2965), .Z(n1979)
         );
  CMX2X4 U4751 ( .A0(\memory[5][37] ), .A1(out_new[37]), .S(N2965), .Z(n1980)
         );
  CMX2X4 U4752 ( .A0(\memory[5][36] ), .A1(out_new[36]), .S(N2965), .Z(n1981)
         );
  CMX2X4 U4753 ( .A0(\memory[5][35] ), .A1(out_new[35]), .S(N2965), .Z(n1982)
         );
  CMX2X4 U4754 ( .A0(\memory[5][34] ), .A1(out_new[34]), .S(N2965), .Z(n1983)
         );
  CMX2X4 U4755 ( .A0(\memory[5][33] ), .A1(out_new[33]), .S(N2965), .Z(n1984)
         );
  CMX2X4 U4756 ( .A0(\memory[5][32] ), .A1(out_new[32]), .S(N2965), .Z(n1985)
         );
  CMX2X4 U4757 ( .A0(\memory[5][31] ), .A1(out_new[31]), .S(N2965), .Z(n1986)
         );
  CMX2X4 U4758 ( .A0(\memory[5][30] ), .A1(out_new[30]), .S(N2965), .Z(n1987)
         );
  CMX2X4 U4759 ( .A0(\memory[5][29] ), .A1(out_new[29]), .S(N2965), .Z(n1988)
         );
  CMX2X4 U4760 ( .A0(\memory[5][28] ), .A1(out_new[28]), .S(N2965), .Z(n1989)
         );
  CMX2X4 U4761 ( .A0(\memory[5][27] ), .A1(out_new[27]), .S(N2965), .Z(n1990)
         );
  CMX2X4 U4762 ( .A0(\memory[5][26] ), .A1(out_new[26]), .S(N2965), .Z(n1991)
         );
  CMX2X4 U4763 ( .A0(\memory[5][25] ), .A1(out_new[25]), .S(N2965), .Z(n1992)
         );
  CMX2X4 U4764 ( .A0(\memory[5][24] ), .A1(out_new[24]), .S(N2965), .Z(n1993)
         );
  CMX2X4 U4765 ( .A0(\memory[5][23] ), .A1(out_new[23]), .S(N2965), .Z(n1994)
         );
  CMX2X4 U4766 ( .A0(\memory[5][22] ), .A1(out_new[22]), .S(N2965), .Z(n1995)
         );
  CMX2X4 U4767 ( .A0(\memory[5][21] ), .A1(out_new[21]), .S(N2965), .Z(n1996)
         );
  CMX2X4 U4768 ( .A0(\memory[5][20] ), .A1(out_new[20]), .S(N2965), .Z(n1997)
         );
  CMX2X4 U4769 ( .A0(\memory[5][19] ), .A1(out_new[19]), .S(N2965), .Z(n1998)
         );
  CMX2X4 U4770 ( .A0(\memory[5][18] ), .A1(out_new[18]), .S(N2965), .Z(n1999)
         );
  CMX2X4 U4771 ( .A0(\memory[5][17] ), .A1(out_new[17]), .S(N2965), .Z(n2000)
         );
  CMX2X4 U4772 ( .A0(\memory[5][16] ), .A1(out_new[16]), .S(N2965), .Z(n2001)
         );
  CMX2X4 U4773 ( .A0(\memory[5][15] ), .A1(out_new[15]), .S(N2965), .Z(n2002)
         );
  CMX2X4 U4774 ( .A0(\memory[5][14] ), .A1(out_new[14]), .S(N2965), .Z(n2003)
         );
  CMX2X4 U4775 ( .A0(\memory[5][13] ), .A1(out_new[13]), .S(N2965), .Z(n2004)
         );
  CMX2X4 U4776 ( .A0(\memory[5][12] ), .A1(out_new[12]), .S(N2965), .Z(n2005)
         );
  CMX2X4 U4777 ( .A0(\memory[5][11] ), .A1(out_new[11]), .S(N2965), .Z(n2006)
         );
  CMX2X4 U4778 ( .A0(\memory[5][10] ), .A1(out_new[10]), .S(N2965), .Z(n2007)
         );
  CMX2X4 U4779 ( .A0(\memory[5][9] ), .A1(out_new[9]), .S(N2965), .Z(n2008) );
  CMX2X4 U4780 ( .A0(\memory[5][8] ), .A1(out_new[8]), .S(N2965), .Z(n2009) );
  CMX2X4 U4781 ( .A0(\memory[5][7] ), .A1(out_new[7]), .S(N2965), .Z(n2010) );
  CMX2X4 U4782 ( .A0(\memory[5][6] ), .A1(out_new[6]), .S(N2965), .Z(n2011) );
  CMX2X4 U4783 ( .A0(\memory[5][5] ), .A1(out_new[5]), .S(N2965), .Z(n2012) );
  CMX2X4 U4784 ( .A0(\memory[5][4] ), .A1(out_new[4]), .S(N2965), .Z(n2013) );
  CMX2X4 U4785 ( .A0(\memory[5][3] ), .A1(out_new[3]), .S(N2965), .Z(n2014) );
  CMX2X4 U4786 ( .A0(\memory[5][2] ), .A1(out_new[2]), .S(N2965), .Z(n2015) );
  CMX2X4 U4787 ( .A0(\memory[5][1] ), .A1(out_new[1]), .S(N2965), .Z(n2016) );
  CMX2X4 U4788 ( .A0(\memory[5][0] ), .A1(out_new[0]), .S(N2965), .Z(n2017) );
  CMX2X2 U4789 ( .A0(\memory[4][63] ), .A1(out_new[63]), .S(N2894), .Z(n2025)
         );
  CMX2X2 U4790 ( .A0(\memory[4][62] ), .A1(out_new[62]), .S(N2894), .Z(n2026)
         );
  CMX2X2 U4791 ( .A0(\memory[4][61] ), .A1(out_new[61]), .S(N2894), .Z(n2027)
         );
  CMX2X2 U4792 ( .A0(\memory[4][60] ), .A1(out_new[60]), .S(N2894), .Z(n2028)
         );
  CMX2X2 U4793 ( .A0(\memory[4][59] ), .A1(out_new[59]), .S(N2894), .Z(n2029)
         );
  CMX2X2 U4794 ( .A0(\memory[4][58] ), .A1(out_new[58]), .S(N2894), .Z(n2030)
         );
  CMX2X2 U4795 ( .A0(\memory[4][57] ), .A1(out_new[57]), .S(N2894), .Z(n2031)
         );
  CMX2X2 U4796 ( .A0(\memory[4][56] ), .A1(out_new[56]), .S(N2894), .Z(n2032)
         );
  CMX2X2 U4797 ( .A0(\memory[4][55] ), .A1(out_new[55]), .S(N2894), .Z(n2033)
         );
  CMX2X2 U4798 ( .A0(\memory[4][54] ), .A1(out_new[54]), .S(N2894), .Z(n2034)
         );
  CMX2X2 U4799 ( .A0(\memory[4][53] ), .A1(out_new[53]), .S(N2894), .Z(n2035)
         );
  CMX2X2 U4800 ( .A0(\memory[4][52] ), .A1(out_new[52]), .S(N2894), .Z(n2036)
         );
  CMX2X2 U4801 ( .A0(\memory[4][51] ), .A1(out_new[51]), .S(N2894), .Z(n2037)
         );
  CMX2X2 U4802 ( .A0(\memory[4][50] ), .A1(out_new[50]), .S(N2894), .Z(n2038)
         );
  CMX2X2 U4803 ( .A0(\memory[4][49] ), .A1(out_new[49]), .S(N2894), .Z(n2039)
         );
  CMX2X2 U4804 ( .A0(\memory[4][48] ), .A1(out_new[48]), .S(N2894), .Z(n2040)
         );
  CMX2X2 U4805 ( .A0(\memory[4][47] ), .A1(out_new[47]), .S(N2894), .Z(n2041)
         );
  CMX2X2 U4806 ( .A0(\memory[4][46] ), .A1(out_new[46]), .S(N2894), .Z(n2042)
         );
  CMX2X2 U4807 ( .A0(\memory[4][45] ), .A1(out_new[45]), .S(N2894), .Z(n2043)
         );
  CMX2X2 U4808 ( .A0(\memory[4][44] ), .A1(out_new[44]), .S(N2894), .Z(n2044)
         );
  CMX2X2 U4809 ( .A0(\memory[4][43] ), .A1(out_new[43]), .S(N2894), .Z(n2045)
         );
  CMX2X2 U4810 ( .A0(\memory[4][42] ), .A1(out_new[42]), .S(N2894), .Z(n2046)
         );
  CMX2X2 U4811 ( .A0(\memory[4][41] ), .A1(out_new[41]), .S(N2894), .Z(n2047)
         );
  CMX2X2 U4812 ( .A0(\memory[4][40] ), .A1(out_new[40]), .S(N2894), .Z(n2048)
         );
  CMX2X2 U4813 ( .A0(\memory[4][39] ), .A1(out_new[39]), .S(N2894), .Z(n2049)
         );
  CMX2X2 U4814 ( .A0(\memory[4][38] ), .A1(out_new[38]), .S(N2894), .Z(n2050)
         );
  CMX2X2 U4815 ( .A0(\memory[4][37] ), .A1(out_new[37]), .S(N2894), .Z(n2051)
         );
  CMX2X2 U4816 ( .A0(\memory[4][36] ), .A1(out_new[36]), .S(N2894), .Z(n2052)
         );
  CMX2X2 U4817 ( .A0(\memory[4][35] ), .A1(out_new[35]), .S(N2894), .Z(n2053)
         );
  CMX2X2 U4818 ( .A0(\memory[4][34] ), .A1(out_new[34]), .S(N2894), .Z(n2054)
         );
  CMX2X2 U4819 ( .A0(\memory[4][33] ), .A1(out_new[33]), .S(N2894), .Z(n2055)
         );
  CMX2X2 U4820 ( .A0(\memory[4][32] ), .A1(out_new[32]), .S(N2894), .Z(n2056)
         );
  CMX2X2 U4821 ( .A0(\memory[4][31] ), .A1(out_new[31]), .S(N2894), .Z(n2057)
         );
  CMX2X2 U4822 ( .A0(\memory[4][30] ), .A1(out_new[30]), .S(N2894), .Z(n2058)
         );
  CMX2X2 U4823 ( .A0(\memory[4][29] ), .A1(out_new[29]), .S(N2894), .Z(n2059)
         );
  CMX2X2 U4824 ( .A0(\memory[4][28] ), .A1(out_new[28]), .S(N2894), .Z(n2060)
         );
  CMX2X2 U4825 ( .A0(\memory[4][27] ), .A1(out_new[27]), .S(N2894), .Z(n2061)
         );
  CMX2X2 U4826 ( .A0(\memory[4][26] ), .A1(out_new[26]), .S(N2894), .Z(n2062)
         );
  CMX2X2 U4827 ( .A0(\memory[4][25] ), .A1(out_new[25]), .S(N2894), .Z(n2063)
         );
  CMX2X2 U4828 ( .A0(\memory[4][24] ), .A1(out_new[24]), .S(N2894), .Z(n2064)
         );
  CMX2X2 U4829 ( .A0(\memory[4][23] ), .A1(out_new[23]), .S(N2894), .Z(n2065)
         );
  CMX2X2 U4830 ( .A0(\memory[4][22] ), .A1(out_new[22]), .S(N2894), .Z(n2066)
         );
  CMX2X2 U4831 ( .A0(\memory[4][21] ), .A1(out_new[21]), .S(N2894), .Z(n2067)
         );
  CMX2X2 U4832 ( .A0(\memory[4][20] ), .A1(out_new[20]), .S(N2894), .Z(n2068)
         );
  CMX2X2 U4833 ( .A0(\memory[4][19] ), .A1(out_new[19]), .S(N2894), .Z(n2069)
         );
  CMX2X2 U4834 ( .A0(\memory[4][18] ), .A1(out_new[18]), .S(N2894), .Z(n2070)
         );
  CMX2X2 U4835 ( .A0(\memory[4][17] ), .A1(out_new[17]), .S(N2894), .Z(n2071)
         );
  CMX2X2 U4836 ( .A0(\memory[4][16] ), .A1(out_new[16]), .S(N2894), .Z(n2072)
         );
  CMX2X2 U4837 ( .A0(\memory[4][15] ), .A1(out_new[15]), .S(N2894), .Z(n2073)
         );
  CMX2X2 U4838 ( .A0(\memory[4][14] ), .A1(out_new[14]), .S(N2894), .Z(n2074)
         );
  CMX2X2 U4839 ( .A0(\memory[4][13] ), .A1(out_new[13]), .S(N2894), .Z(n2075)
         );
  CMX2X2 U4840 ( .A0(\memory[4][12] ), .A1(out_new[12]), .S(N2894), .Z(n2076)
         );
  CMX2X2 U4841 ( .A0(\memory[4][11] ), .A1(out_new[11]), .S(N2894), .Z(n2077)
         );
  CMX2X2 U4842 ( .A0(\memory[4][10] ), .A1(out_new[10]), .S(N2894), .Z(n2078)
         );
  CMX2X2 U4843 ( .A0(\memory[4][9] ), .A1(out_new[9]), .S(N2894), .Z(n2079) );
  CMX2X2 U4844 ( .A0(\memory[4][8] ), .A1(out_new[8]), .S(N2894), .Z(n2080) );
  CMX2X2 U4845 ( .A0(\memory[4][7] ), .A1(out_new[7]), .S(N2894), .Z(n2081) );
  CMX2X2 U4846 ( .A0(\memory[4][6] ), .A1(out_new[6]), .S(N2894), .Z(n2082) );
  CMX2X2 U4847 ( .A0(\memory[4][5] ), .A1(out_new[5]), .S(N2894), .Z(n2083) );
  CMX2X2 U4848 ( .A0(\memory[4][4] ), .A1(out_new[4]), .S(N2894), .Z(n2084) );
  CMX2X2 U4849 ( .A0(\memory[4][3] ), .A1(out_new[3]), .S(N2894), .Z(n2085) );
  CMX2X2 U4850 ( .A0(\memory[4][2] ), .A1(out_new[2]), .S(N2894), .Z(n2086) );
  CMX2X2 U4851 ( .A0(\memory[4][1] ), .A1(out_new[1]), .S(N2894), .Z(n2087) );
  CMX2X2 U4852 ( .A0(\memory[4][0] ), .A1(out_new[0]), .S(N2894), .Z(n2088) );
  CMX2X2 U4853 ( .A0(\memory[3][63] ), .A1(out_new[63]), .S(N2823), .Z(n2096)
         );
  CMX2X2 U4854 ( .A0(\memory[3][62] ), .A1(out_new[62]), .S(N2823), .Z(n2097)
         );
  CMX2X2 U4855 ( .A0(\memory[3][61] ), .A1(out_new[61]), .S(N2823), .Z(n2098)
         );
  CMX2X2 U4856 ( .A0(\memory[3][60] ), .A1(out_new[60]), .S(N2823), .Z(n2099)
         );
  CMX2X2 U4857 ( .A0(\memory[3][59] ), .A1(out_new[59]), .S(N2823), .Z(n2100)
         );
  CMX2X2 U4858 ( .A0(\memory[3][58] ), .A1(out_new[58]), .S(N2823), .Z(n2101)
         );
  CMX2X2 U4859 ( .A0(\memory[3][57] ), .A1(out_new[57]), .S(N2823), .Z(n2102)
         );
  CMX2X2 U4860 ( .A0(\memory[3][56] ), .A1(out_new[56]), .S(N2823), .Z(n2103)
         );
  CMX2X2 U4861 ( .A0(\memory[3][55] ), .A1(out_new[55]), .S(N2823), .Z(n2104)
         );
  CMX2X2 U4862 ( .A0(\memory[3][54] ), .A1(out_new[54]), .S(N2823), .Z(n2105)
         );
  CMX2X2 U4863 ( .A0(\memory[3][53] ), .A1(out_new[53]), .S(N2823), .Z(n2106)
         );
  CMX2X2 U4864 ( .A0(\memory[3][52] ), .A1(out_new[52]), .S(N2823), .Z(n2107)
         );
  CMX2X2 U4865 ( .A0(\memory[3][51] ), .A1(out_new[51]), .S(N2823), .Z(n2108)
         );
  CMX2X2 U4866 ( .A0(\memory[3][50] ), .A1(out_new[50]), .S(N2823), .Z(n2109)
         );
  CMX2X2 U4867 ( .A0(\memory[3][49] ), .A1(out_new[49]), .S(N2823), .Z(n2110)
         );
  CMX2X2 U4868 ( .A0(\memory[3][48] ), .A1(out_new[48]), .S(N2823), .Z(n2111)
         );
  CMX2X2 U4869 ( .A0(\memory[3][47] ), .A1(out_new[47]), .S(N2823), .Z(n2112)
         );
  CMX2X2 U4870 ( .A0(\memory[3][46] ), .A1(out_new[46]), .S(N2823), .Z(n2113)
         );
  CMX2X2 U4871 ( .A0(\memory[3][45] ), .A1(out_new[45]), .S(N2823), .Z(n2114)
         );
  CMX2X2 U4872 ( .A0(\memory[3][44] ), .A1(out_new[44]), .S(N2823), .Z(n2115)
         );
  CMX2X2 U4873 ( .A0(\memory[3][43] ), .A1(out_new[43]), .S(N2823), .Z(n2116)
         );
  CMX2X2 U4874 ( .A0(\memory[3][42] ), .A1(out_new[42]), .S(N2823), .Z(n2117)
         );
  CMX2X2 U4875 ( .A0(\memory[3][41] ), .A1(out_new[41]), .S(N2823), .Z(n2118)
         );
  CMX2X2 U4876 ( .A0(\memory[3][40] ), .A1(out_new[40]), .S(N2823), .Z(n2119)
         );
  CMX2X2 U4877 ( .A0(\memory[3][39] ), .A1(out_new[39]), .S(N2823), .Z(n2120)
         );
  CMX2X2 U4878 ( .A0(\memory[3][38] ), .A1(out_new[38]), .S(N2823), .Z(n2121)
         );
  CMX2X2 U4879 ( .A0(\memory[3][37] ), .A1(out_new[37]), .S(N2823), .Z(n2122)
         );
  CMX2X2 U4880 ( .A0(\memory[3][36] ), .A1(out_new[36]), .S(N2823), .Z(n2123)
         );
  CMX2X2 U4881 ( .A0(\memory[3][35] ), .A1(out_new[35]), .S(N2823), .Z(n2124)
         );
  CMX2X2 U4882 ( .A0(\memory[3][34] ), .A1(out_new[34]), .S(N2823), .Z(n2125)
         );
  CMX2X2 U4883 ( .A0(\memory[3][33] ), .A1(out_new[33]), .S(N2823), .Z(n2126)
         );
  CMX2X2 U4884 ( .A0(\memory[3][32] ), .A1(out_new[32]), .S(N2823), .Z(n2127)
         );
  CMX2X2 U4885 ( .A0(\memory[3][31] ), .A1(out_new[31]), .S(N2823), .Z(n2128)
         );
  CMX2X2 U4886 ( .A0(\memory[3][30] ), .A1(out_new[30]), .S(N2823), .Z(n2129)
         );
  CMX2X2 U4887 ( .A0(\memory[3][29] ), .A1(out_new[29]), .S(N2823), .Z(n2130)
         );
  CMX2X2 U4888 ( .A0(\memory[3][28] ), .A1(out_new[28]), .S(N2823), .Z(n2131)
         );
  CMX2X2 U4889 ( .A0(\memory[3][27] ), .A1(out_new[27]), .S(N2823), .Z(n2132)
         );
  CMX2X2 U4890 ( .A0(\memory[3][26] ), .A1(out_new[26]), .S(N2823), .Z(n2133)
         );
  CMX2X2 U4891 ( .A0(\memory[3][25] ), .A1(out_new[25]), .S(N2823), .Z(n2134)
         );
  CMX2X2 U4892 ( .A0(\memory[3][24] ), .A1(out_new[24]), .S(N2823), .Z(n2135)
         );
  CMX2X2 U4893 ( .A0(\memory[3][23] ), .A1(out_new[23]), .S(N2823), .Z(n2136)
         );
  CMX2X2 U4894 ( .A0(\memory[3][22] ), .A1(out_new[22]), .S(N2823), .Z(n2137)
         );
  CMX2X2 U4895 ( .A0(\memory[3][21] ), .A1(out_new[21]), .S(N2823), .Z(n2138)
         );
  CMX2X2 U4896 ( .A0(\memory[3][20] ), .A1(out_new[20]), .S(N2823), .Z(n2139)
         );
  CMX2X2 U4897 ( .A0(\memory[3][19] ), .A1(out_new[19]), .S(N2823), .Z(n2140)
         );
  CMX2X2 U4898 ( .A0(\memory[3][18] ), .A1(out_new[18]), .S(N2823), .Z(n2141)
         );
  CMX2X2 U4899 ( .A0(\memory[3][17] ), .A1(out_new[17]), .S(N2823), .Z(n2142)
         );
  CMX2X2 U4900 ( .A0(\memory[3][16] ), .A1(out_new[16]), .S(N2823), .Z(n2143)
         );
  CMX2X2 U4901 ( .A0(\memory[3][15] ), .A1(out_new[15]), .S(N2823), .Z(n2144)
         );
  CMX2X2 U4902 ( .A0(\memory[3][14] ), .A1(out_new[14]), .S(N2823), .Z(n2145)
         );
  CMX2X2 U4903 ( .A0(\memory[3][13] ), .A1(out_new[13]), .S(N2823), .Z(n2146)
         );
  CMX2X2 U4904 ( .A0(\memory[3][12] ), .A1(out_new[12]), .S(N2823), .Z(n2147)
         );
  CMX2X2 U4905 ( .A0(\memory[3][11] ), .A1(out_new[11]), .S(N2823), .Z(n2148)
         );
  CMX2X2 U4906 ( .A0(\memory[3][10] ), .A1(out_new[10]), .S(N2823), .Z(n2149)
         );
  CMX2X2 U4907 ( .A0(\memory[3][9] ), .A1(out_new[9]), .S(N2823), .Z(n2150) );
  CMX2X2 U4908 ( .A0(\memory[3][8] ), .A1(out_new[8]), .S(N2823), .Z(n2151) );
  CMX2X2 U4909 ( .A0(\memory[3][7] ), .A1(out_new[7]), .S(N2823), .Z(n2152) );
  CMX2X2 U4910 ( .A0(\memory[3][6] ), .A1(out_new[6]), .S(N2823), .Z(n2153) );
  CMX2X2 U4911 ( .A0(\memory[3][5] ), .A1(out_new[5]), .S(N2823), .Z(n2154) );
  CMX2X2 U4912 ( .A0(\memory[3][4] ), .A1(out_new[4]), .S(N2823), .Z(n2155) );
  CMX2X2 U4913 ( .A0(\memory[3][3] ), .A1(out_new[3]), .S(N2823), .Z(n2156) );
  CMX2X2 U4914 ( .A0(\memory[3][2] ), .A1(out_new[2]), .S(N2823), .Z(n2157) );
  CMX2X2 U4915 ( .A0(\memory[3][1] ), .A1(out_new[1]), .S(N2823), .Z(n2158) );
  CMX2X2 U4916 ( .A0(\memory[3][0] ), .A1(out_new[0]), .S(N2823), .Z(n2159) );
  CMX2X2 U4917 ( .A0(\memory[2][63] ), .A1(out_new[63]), .S(n2603), .Z(n2167)
         );
  CMX2X2 U4918 ( .A0(\memory[2][62] ), .A1(out_new[62]), .S(n2603), .Z(n2168)
         );
  CMX2X2 U4919 ( .A0(\memory[2][61] ), .A1(out_new[61]), .S(n2603), .Z(n2169)
         );
  CMX2X2 U4920 ( .A0(\memory[2][60] ), .A1(out_new[60]), .S(n2603), .Z(n2170)
         );
  CMX2X2 U4921 ( .A0(\memory[2][59] ), .A1(out_new[59]), .S(n2603), .Z(n2171)
         );
  CMX2X2 U4922 ( .A0(\memory[2][58] ), .A1(out_new[58]), .S(n2603), .Z(n2172)
         );
  CMX2X2 U4923 ( .A0(\memory[2][57] ), .A1(out_new[57]), .S(n2603), .Z(n2173)
         );
  CMX2X2 U4924 ( .A0(\memory[2][56] ), .A1(out_new[56]), .S(n2603), .Z(n2174)
         );
  CMX2X2 U4925 ( .A0(\memory[2][55] ), .A1(out_new[55]), .S(n2603), .Z(n2175)
         );
  CMX2X2 U4926 ( .A0(\memory[2][54] ), .A1(out_new[54]), .S(n2603), .Z(n2176)
         );
  CMX2X2 U4927 ( .A0(\memory[2][53] ), .A1(out_new[53]), .S(n2603), .Z(n2177)
         );
  CMX2X2 U4928 ( .A0(\memory[2][52] ), .A1(out_new[52]), .S(n2603), .Z(n2178)
         );
  CMX2X2 U4929 ( .A0(\memory[2][51] ), .A1(out_new[51]), .S(n2603), .Z(n2179)
         );
  CMX2X2 U4930 ( .A0(\memory[2][50] ), .A1(out_new[50]), .S(n2603), .Z(n2180)
         );
  CMX2X2 U4931 ( .A0(\memory[2][49] ), .A1(out_new[49]), .S(n2603), .Z(n2181)
         );
  CMX2X2 U4932 ( .A0(\memory[2][48] ), .A1(out_new[48]), .S(n2603), .Z(n2182)
         );
  CMX2X2 U4933 ( .A0(\memory[2][47] ), .A1(out_new[47]), .S(n2603), .Z(n2183)
         );
  CMX2X2 U4934 ( .A0(\memory[2][46] ), .A1(out_new[46]), .S(n2603), .Z(n2184)
         );
  CMX2X2 U4935 ( .A0(\memory[2][45] ), .A1(out_new[45]), .S(n2603), .Z(n2185)
         );
  CMX2X2 U4936 ( .A0(\memory[2][44] ), .A1(out_new[44]), .S(n2603), .Z(n2186)
         );
  CMX2X2 U4937 ( .A0(\memory[2][43] ), .A1(out_new[43]), .S(n2603), .Z(n2187)
         );
  CMX2X2 U4938 ( .A0(\memory[2][42] ), .A1(out_new[42]), .S(n2603), .Z(n2188)
         );
  CMX2X2 U4939 ( .A0(\memory[2][41] ), .A1(out_new[41]), .S(n2603), .Z(n2189)
         );
  CMX2X2 U4940 ( .A0(\memory[2][40] ), .A1(out_new[40]), .S(n2603), .Z(n2190)
         );
  CMX2X2 U4941 ( .A0(\memory[2][39] ), .A1(out_new[39]), .S(n2603), .Z(n2191)
         );
  CMX2X2 U4942 ( .A0(\memory[2][38] ), .A1(out_new[38]), .S(n2603), .Z(n2192)
         );
  CMX2X2 U4943 ( .A0(\memory[2][37] ), .A1(out_new[37]), .S(n2603), .Z(n2193)
         );
  CMX2X2 U4944 ( .A0(\memory[2][36] ), .A1(out_new[36]), .S(n2603), .Z(n2194)
         );
  CMX2X2 U4945 ( .A0(\memory[2][35] ), .A1(out_new[35]), .S(n2603), .Z(n2195)
         );
  CMX2X2 U4946 ( .A0(\memory[2][34] ), .A1(out_new[34]), .S(n2603), .Z(n2196)
         );
  CMX2X2 U4947 ( .A0(\memory[2][33] ), .A1(out_new[33]), .S(n2603), .Z(n2197)
         );
  CMX2X2 U4948 ( .A0(\memory[2][32] ), .A1(out_new[32]), .S(n2603), .Z(n2198)
         );
  CMX2X2 U4949 ( .A0(\memory[2][31] ), .A1(out_new[31]), .S(n2603), .Z(n2199)
         );
  CMX2X2 U4950 ( .A0(\memory[2][30] ), .A1(out_new[30]), .S(n2603), .Z(n2200)
         );
  CMX2X2 U4951 ( .A0(\memory[2][29] ), .A1(out_new[29]), .S(n2603), .Z(n2201)
         );
  CMX2X2 U4952 ( .A0(\memory[2][28] ), .A1(out_new[28]), .S(n2603), .Z(n2202)
         );
  CMX2X2 U4953 ( .A0(\memory[2][27] ), .A1(out_new[27]), .S(n2603), .Z(n2203)
         );
  CMX2X2 U4954 ( .A0(\memory[2][26] ), .A1(out_new[26]), .S(n2603), .Z(n2204)
         );
  CMX2X2 U4955 ( .A0(\memory[2][25] ), .A1(out_new[25]), .S(n2603), .Z(n2205)
         );
  CMX2X2 U4956 ( .A0(\memory[2][24] ), .A1(out_new[24]), .S(n2603), .Z(n2206)
         );
  CMX2X2 U4957 ( .A0(\memory[2][23] ), .A1(out_new[23]), .S(n2603), .Z(n2207)
         );
  CMX2X2 U4958 ( .A0(\memory[2][22] ), .A1(out_new[22]), .S(n2603), .Z(n2208)
         );
  CMX2X2 U4959 ( .A0(\memory[2][21] ), .A1(out_new[21]), .S(n2603), .Z(n2209)
         );
  CMX2X2 U4960 ( .A0(\memory[2][20] ), .A1(out_new[20]), .S(n2603), .Z(n2210)
         );
  CMX2X2 U4961 ( .A0(\memory[2][19] ), .A1(out_new[19]), .S(n2603), .Z(n2211)
         );
  CMX2X2 U4962 ( .A0(\memory[2][18] ), .A1(out_new[18]), .S(n2603), .Z(n2212)
         );
  CMX2X2 U4963 ( .A0(\memory[2][17] ), .A1(out_new[17]), .S(n2603), .Z(n2213)
         );
  CMX2X2 U4964 ( .A0(\memory[2][16] ), .A1(out_new[16]), .S(n2603), .Z(n2214)
         );
  CMX2X2 U4965 ( .A0(\memory[2][15] ), .A1(out_new[15]), .S(n2603), .Z(n2215)
         );
  CMX2X2 U4966 ( .A0(\memory[2][14] ), .A1(out_new[14]), .S(n2603), .Z(n2216)
         );
  CMX2X2 U4967 ( .A0(\memory[2][13] ), .A1(out_new[13]), .S(n2603), .Z(n2217)
         );
  CMX2X2 U4968 ( .A0(\memory[2][12] ), .A1(out_new[12]), .S(n2603), .Z(n2218)
         );
  CMX2X2 U4969 ( .A0(\memory[2][11] ), .A1(out_new[11]), .S(n2603), .Z(n2219)
         );
  CMX2X2 U4970 ( .A0(\memory[2][10] ), .A1(out_new[10]), .S(n2603), .Z(n2220)
         );
  CMX2X2 U4971 ( .A0(\memory[2][9] ), .A1(out_new[9]), .S(n2603), .Z(n2221) );
  CMX2X2 U4972 ( .A0(\memory[2][8] ), .A1(out_new[8]), .S(n2603), .Z(n2222) );
  CMX2X2 U4973 ( .A0(\memory[2][7] ), .A1(out_new[7]), .S(n2603), .Z(n2223) );
  CMX2X2 U4974 ( .A0(\memory[2][6] ), .A1(out_new[6]), .S(n2603), .Z(n2224) );
  CMX2X2 U4975 ( .A0(\memory[2][5] ), .A1(out_new[5]), .S(n2603), .Z(n2225) );
  CMX2X2 U4976 ( .A0(\memory[2][4] ), .A1(out_new[4]), .S(n2603), .Z(n2226) );
  CMX2X2 U4977 ( .A0(\memory[2][3] ), .A1(out_new[3]), .S(n2603), .Z(n2227) );
  CMX2X2 U4978 ( .A0(\memory[2][2] ), .A1(out_new[2]), .S(n2603), .Z(n2228) );
  CMX2X2 U4979 ( .A0(\memory[2][1] ), .A1(out_new[1]), .S(n2603), .Z(n2229) );
  CMX2X2 U4980 ( .A0(\memory[2][0] ), .A1(out_new[0]), .S(n2603), .Z(n2230) );
  CMX2X2 U4981 ( .A0(\memory[1][63] ), .A1(out_new[63]), .S(n2601), .Z(n2238)
         );
  CMX2X2 U4982 ( .A0(\memory[1][62] ), .A1(out_new[62]), .S(n2601), .Z(n2239)
         );
  CMX2X2 U4983 ( .A0(\memory[1][61] ), .A1(out_new[61]), .S(n2601), .Z(n2240)
         );
  CMX2X2 U4984 ( .A0(\memory[1][60] ), .A1(out_new[60]), .S(n2601), .Z(n2241)
         );
  CMX2X2 U4985 ( .A0(\memory[1][59] ), .A1(out_new[59]), .S(n2601), .Z(n2242)
         );
  CMX2X2 U4986 ( .A0(\memory[1][58] ), .A1(out_new[58]), .S(n2601), .Z(n2243)
         );
  CMX2X2 U4987 ( .A0(\memory[1][57] ), .A1(out_new[57]), .S(n2601), .Z(n2244)
         );
  CMX2X2 U4988 ( .A0(\memory[1][56] ), .A1(out_new[56]), .S(n2601), .Z(n2245)
         );
  CMX2X2 U4989 ( .A0(\memory[1][55] ), .A1(out_new[55]), .S(n2601), .Z(n2246)
         );
  CMX2X2 U4990 ( .A0(\memory[1][54] ), .A1(out_new[54]), .S(n2601), .Z(n2247)
         );
  CMX2X2 U4991 ( .A0(\memory[1][53] ), .A1(out_new[53]), .S(n2601), .Z(n2248)
         );
  CMX2X2 U4992 ( .A0(\memory[1][52] ), .A1(out_new[52]), .S(n2601), .Z(n2249)
         );
  CMX2X2 U4993 ( .A0(\memory[1][51] ), .A1(out_new[51]), .S(n2601), .Z(n2250)
         );
  CMX2X2 U4994 ( .A0(\memory[1][50] ), .A1(out_new[50]), .S(n2601), .Z(n2251)
         );
  CMX2X2 U4995 ( .A0(\memory[1][49] ), .A1(out_new[49]), .S(n2601), .Z(n2252)
         );
  CMX2X2 U4996 ( .A0(\memory[1][48] ), .A1(out_new[48]), .S(n2601), .Z(n2253)
         );
  CMX2X2 U4997 ( .A0(\memory[1][47] ), .A1(out_new[47]), .S(n2601), .Z(n2254)
         );
  CMX2X2 U4998 ( .A0(\memory[1][46] ), .A1(out_new[46]), .S(n2601), .Z(n2255)
         );
  CMX2X2 U4999 ( .A0(\memory[1][45] ), .A1(out_new[45]), .S(n2601), .Z(n2256)
         );
  CMX2X2 U5000 ( .A0(\memory[1][44] ), .A1(out_new[44]), .S(n2601), .Z(n2257)
         );
  CMX2X2 U5001 ( .A0(\memory[1][43] ), .A1(out_new[43]), .S(n2601), .Z(n2258)
         );
  CMX2X2 U5002 ( .A0(\memory[1][42] ), .A1(out_new[42]), .S(n2601), .Z(n2259)
         );
  CMX2X2 U5003 ( .A0(\memory[1][41] ), .A1(out_new[41]), .S(n2601), .Z(n2260)
         );
  CMX2X2 U5004 ( .A0(\memory[1][40] ), .A1(out_new[40]), .S(n2601), .Z(n2261)
         );
  CMX2X2 U5005 ( .A0(\memory[1][39] ), .A1(out_new[39]), .S(n2601), .Z(n2262)
         );
  CMX2X2 U5006 ( .A0(\memory[1][38] ), .A1(out_new[38]), .S(n2601), .Z(n2263)
         );
  CMX2X2 U5007 ( .A0(\memory[1][37] ), .A1(out_new[37]), .S(n2601), .Z(n2264)
         );
  CMX2X2 U5008 ( .A0(\memory[1][36] ), .A1(out_new[36]), .S(n2601), .Z(n2265)
         );
  CMX2X2 U5009 ( .A0(\memory[1][35] ), .A1(out_new[35]), .S(n2601), .Z(n2266)
         );
  CMX2X2 U5010 ( .A0(\memory[1][34] ), .A1(out_new[34]), .S(n2601), .Z(n2267)
         );
  CMX2X2 U5011 ( .A0(\memory[1][33] ), .A1(out_new[33]), .S(n2601), .Z(n2268)
         );
  CMX2X2 U5012 ( .A0(\memory[1][32] ), .A1(out_new[32]), .S(n2601), .Z(n2269)
         );
  CMX2X2 U5013 ( .A0(\memory[1][31] ), .A1(out_new[31]), .S(n2601), .Z(n2270)
         );
  CMX2X2 U5014 ( .A0(\memory[1][30] ), .A1(out_new[30]), .S(n2601), .Z(n2271)
         );
  CMX2X2 U5015 ( .A0(\memory[1][29] ), .A1(out_new[29]), .S(n2601), .Z(n2272)
         );
  CMX2X2 U5016 ( .A0(\memory[1][28] ), .A1(out_new[28]), .S(n2601), .Z(n2273)
         );
  CMX2X2 U5017 ( .A0(\memory[1][27] ), .A1(out_new[27]), .S(n2601), .Z(n2274)
         );
  CMX2X2 U5018 ( .A0(\memory[1][26] ), .A1(out_new[26]), .S(n2601), .Z(n2275)
         );
  CMX2X2 U5019 ( .A0(\memory[1][25] ), .A1(out_new[25]), .S(n2601), .Z(n2276)
         );
  CMX2X2 U5020 ( .A0(\memory[1][24] ), .A1(out_new[24]), .S(n2601), .Z(n2277)
         );
  CMX2X2 U5021 ( .A0(\memory[1][23] ), .A1(out_new[23]), .S(n2601), .Z(n2278)
         );
  CMX2X2 U5022 ( .A0(\memory[1][22] ), .A1(out_new[22]), .S(n2601), .Z(n2279)
         );
  CMX2X2 U5023 ( .A0(\memory[1][21] ), .A1(out_new[21]), .S(n2601), .Z(n2280)
         );
  CMX2X2 U5024 ( .A0(\memory[1][20] ), .A1(out_new[20]), .S(n2601), .Z(n2281)
         );
  CMX2X2 U5025 ( .A0(\memory[1][19] ), .A1(out_new[19]), .S(n2601), .Z(n2282)
         );
  CMX2X2 U5026 ( .A0(\memory[1][18] ), .A1(out_new[18]), .S(n2601), .Z(n2283)
         );
  CMX2X2 U5027 ( .A0(\memory[1][17] ), .A1(out_new[17]), .S(n2601), .Z(n2284)
         );
  CMX2X2 U5028 ( .A0(\memory[1][16] ), .A1(out_new[16]), .S(n2601), .Z(n2285)
         );
  CMX2X2 U5029 ( .A0(\memory[1][15] ), .A1(out_new[15]), .S(n2601), .Z(n2286)
         );
  CMX2X2 U5030 ( .A0(\memory[1][14] ), .A1(out_new[14]), .S(n2601), .Z(n2287)
         );
  CMX2X2 U5031 ( .A0(\memory[1][13] ), .A1(out_new[13]), .S(n2601), .Z(n2288)
         );
  CMX2X2 U5032 ( .A0(\memory[1][12] ), .A1(out_new[12]), .S(n2601), .Z(n2289)
         );
  CMX2X2 U5033 ( .A0(\memory[1][11] ), .A1(out_new[11]), .S(n2601), .Z(n2290)
         );
  CMX2X2 U5034 ( .A0(\memory[1][10] ), .A1(out_new[10]), .S(n2601), .Z(n2291)
         );
  CMX2X2 U5035 ( .A0(\memory[1][9] ), .A1(out_new[9]), .S(n2601), .Z(n2292) );
  CMX2X2 U5036 ( .A0(\memory[1][8] ), .A1(out_new[8]), .S(n2601), .Z(n2293) );
  CMX2X2 U5037 ( .A0(\memory[1][7] ), .A1(out_new[7]), .S(n2601), .Z(n2294) );
  CMX2X2 U5038 ( .A0(\memory[1][6] ), .A1(out_new[6]), .S(n2601), .Z(n2295) );
  CMX2X2 U5039 ( .A0(\memory[1][5] ), .A1(out_new[5]), .S(n2601), .Z(n2296) );
  CMX2X2 U5040 ( .A0(\memory[1][4] ), .A1(out_new[4]), .S(n2601), .Z(n2297) );
  CMX2X2 U5041 ( .A0(\memory[1][3] ), .A1(out_new[3]), .S(n2601), .Z(n2298) );
  CMX2X2 U5042 ( .A0(\memory[1][2] ), .A1(out_new[2]), .S(n2601), .Z(n2299) );
  CMX2X2 U5043 ( .A0(\memory[1][1] ), .A1(out_new[1]), .S(n2601), .Z(n2300) );
  CMX2X2 U5044 ( .A0(\memory[1][0] ), .A1(out_new[0]), .S(n2601), .Z(n2301) );
  CMX2X2 U5045 ( .A0(\memory[0][63] ), .A1(out_new[63]), .S(n2605), .Z(n2309)
         );
  CMX2X2 U5046 ( .A0(\memory[0][62] ), .A1(out_new[62]), .S(n2605), .Z(n2310)
         );
  CMX2X2 U5047 ( .A0(\memory[0][61] ), .A1(out_new[61]), .S(n2605), .Z(n2311)
         );
  CMX2X2 U5048 ( .A0(\memory[0][60] ), .A1(out_new[60]), .S(n2605), .Z(n2312)
         );
  CMX2X2 U5049 ( .A0(\memory[0][59] ), .A1(out_new[59]), .S(n2605), .Z(n2313)
         );
  CMX2X2 U5050 ( .A0(\memory[0][58] ), .A1(out_new[58]), .S(n2605), .Z(n2314)
         );
  CMX2X2 U5051 ( .A0(\memory[0][57] ), .A1(out_new[57]), .S(n2605), .Z(n2315)
         );
  CMX2X2 U5052 ( .A0(\memory[0][56] ), .A1(out_new[56]), .S(n2605), .Z(n2316)
         );
  CMX2X2 U5053 ( .A0(\memory[0][55] ), .A1(out_new[55]), .S(n2605), .Z(n2317)
         );
  CMX2X2 U5054 ( .A0(\memory[0][54] ), .A1(out_new[54]), .S(n2605), .Z(n2318)
         );
  CMX2X2 U5055 ( .A0(\memory[0][53] ), .A1(out_new[53]), .S(n2605), .Z(n2319)
         );
  CMX2X2 U5056 ( .A0(\memory[0][52] ), .A1(out_new[52]), .S(n2605), .Z(n2320)
         );
  CMX2X2 U5057 ( .A0(\memory[0][51] ), .A1(out_new[51]), .S(n2605), .Z(n2321)
         );
  CMX2X2 U5058 ( .A0(\memory[0][50] ), .A1(out_new[50]), .S(n2605), .Z(n2322)
         );
  CMX2X2 U5059 ( .A0(\memory[0][49] ), .A1(out_new[49]), .S(n2605), .Z(n2323)
         );
  CMX2X2 U5060 ( .A0(\memory[0][48] ), .A1(out_new[48]), .S(n2605), .Z(n2324)
         );
  CMX2X2 U5061 ( .A0(\memory[0][47] ), .A1(out_new[47]), .S(n2605), .Z(n2325)
         );
  CMX2X2 U5062 ( .A0(\memory[0][46] ), .A1(out_new[46]), .S(n2605), .Z(n2326)
         );
  CMX2X2 U5063 ( .A0(\memory[0][45] ), .A1(out_new[45]), .S(n2605), .Z(n2327)
         );
  CMX2X2 U5064 ( .A0(\memory[0][44] ), .A1(out_new[44]), .S(n2605), .Z(n2328)
         );
  CMX2X2 U5065 ( .A0(\memory[0][43] ), .A1(out_new[43]), .S(n2605), .Z(n2329)
         );
  CMX2X2 U5066 ( .A0(\memory[0][42] ), .A1(out_new[42]), .S(n2605), .Z(n2330)
         );
  CMX2X2 U5067 ( .A0(\memory[0][41] ), .A1(out_new[41]), .S(n2605), .Z(n2331)
         );
  CMX2X2 U5068 ( .A0(\memory[0][40] ), .A1(out_new[40]), .S(n2605), .Z(n2332)
         );
  CMX2X2 U5069 ( .A0(\memory[0][39] ), .A1(out_new[39]), .S(n2605), .Z(n2333)
         );
  CMX2X2 U5070 ( .A0(\memory[0][38] ), .A1(out_new[38]), .S(n2605), .Z(n2334)
         );
  CMX2X2 U5071 ( .A0(\memory[0][37] ), .A1(out_new[37]), .S(n2605), .Z(n2335)
         );
  CMX2X2 U5072 ( .A0(\memory[0][36] ), .A1(out_new[36]), .S(n2605), .Z(n2336)
         );
  CMX2X2 U5073 ( .A0(\memory[0][35] ), .A1(out_new[35]), .S(n2605), .Z(n2337)
         );
  CMX2X2 U5074 ( .A0(\memory[0][34] ), .A1(out_new[34]), .S(n2605), .Z(n2338)
         );
  CMX2X2 U5075 ( .A0(\memory[0][33] ), .A1(out_new[33]), .S(n2605), .Z(n2339)
         );
  CMX2X2 U5076 ( .A0(\memory[0][32] ), .A1(out_new[32]), .S(n2605), .Z(n2340)
         );
  CMX2X2 U5077 ( .A0(\memory[0][31] ), .A1(out_new[31]), .S(n2605), .Z(n2341)
         );
  CMX2X2 U5078 ( .A0(\memory[0][30] ), .A1(out_new[30]), .S(n2605), .Z(n2342)
         );
  CMX2X2 U5079 ( .A0(\memory[0][29] ), .A1(out_new[29]), .S(n2605), .Z(n2343)
         );
  CMX2X2 U5080 ( .A0(\memory[0][28] ), .A1(out_new[28]), .S(n2605), .Z(n2344)
         );
  CMX2X2 U5081 ( .A0(\memory[0][27] ), .A1(out_new[27]), .S(n2605), .Z(n2345)
         );
  CMX2X2 U5082 ( .A0(\memory[0][26] ), .A1(out_new[26]), .S(n2605), .Z(n2346)
         );
  CMX2X2 U5083 ( .A0(\memory[0][25] ), .A1(out_new[25]), .S(n2605), .Z(n2347)
         );
  CMX2X2 U5084 ( .A0(\memory[0][24] ), .A1(out_new[24]), .S(n2605), .Z(n2348)
         );
  CMX2X2 U5085 ( .A0(\memory[0][23] ), .A1(out_new[23]), .S(n2605), .Z(n2349)
         );
  CMX2X2 U5086 ( .A0(\memory[0][22] ), .A1(out_new[22]), .S(n2605), .Z(n2350)
         );
  CMX2X2 U5087 ( .A0(\memory[0][21] ), .A1(out_new[21]), .S(n2605), .Z(n2351)
         );
  CMX2X2 U5088 ( .A0(\memory[0][20] ), .A1(out_new[20]), .S(n2605), .Z(n2352)
         );
  CMX2X2 U5089 ( .A0(\memory[0][19] ), .A1(out_new[19]), .S(n2605), .Z(n2353)
         );
  CMX2X2 U5090 ( .A0(\memory[0][18] ), .A1(out_new[18]), .S(n2605), .Z(n2354)
         );
  CMX2X2 U5091 ( .A0(\memory[0][17] ), .A1(out_new[17]), .S(n2605), .Z(n2355)
         );
  CMX2X2 U5092 ( .A0(\memory[0][16] ), .A1(out_new[16]), .S(n2605), .Z(n2356)
         );
  CMX2X2 U5093 ( .A0(\memory[0][15] ), .A1(out_new[15]), .S(n2605), .Z(n2357)
         );
  CMX2X2 U5094 ( .A0(\memory[0][14] ), .A1(out_new[14]), .S(n2605), .Z(n2358)
         );
  CMX2X2 U5095 ( .A0(\memory[0][13] ), .A1(out_new[13]), .S(n2605), .Z(n2359)
         );
  CMX2X2 U5096 ( .A0(\memory[0][12] ), .A1(out_new[12]), .S(n2605), .Z(n2360)
         );
  CMX2X2 U5097 ( .A0(\memory[0][11] ), .A1(out_new[11]), .S(n2605), .Z(n2361)
         );
  CMX2X2 U5098 ( .A0(\memory[0][10] ), .A1(out_new[10]), .S(n2605), .Z(n2362)
         );
  CMX2X2 U5099 ( .A0(\memory[0][9] ), .A1(out_new[9]), .S(n2605), .Z(n2363) );
  CMX2X2 U5100 ( .A0(\memory[0][8] ), .A1(out_new[8]), .S(n2605), .Z(n2364) );
  CMX2X2 U5101 ( .A0(\memory[0][7] ), .A1(out_new[7]), .S(n2605), .Z(n2365) );
  CMX2X2 U5102 ( .A0(\memory[0][6] ), .A1(out_new[6]), .S(n2605), .Z(n2366) );
  CMX2X2 U5103 ( .A0(\memory[0][5] ), .A1(out_new[5]), .S(n2605), .Z(n2367) );
  CMX2X2 U5104 ( .A0(\memory[0][4] ), .A1(out_new[4]), .S(n2605), .Z(n2368) );
  CMX2X2 U5105 ( .A0(\memory[0][3] ), .A1(out_new[3]), .S(n2605), .Z(n2369) );
  CMX2X2 U5106 ( .A0(\memory[0][2] ), .A1(out_new[2]), .S(n2605), .Z(n2370) );
  CMX2X2 U5107 ( .A0(\memory[0][1] ), .A1(out_new[1]), .S(n2605), .Z(n2371) );
  CMX2X2 U5108 ( .A0(\memory[0][0] ), .A1(out_new[0]), .S(n2605), .Z(n2372) );
  CND2X2 U5109 ( .A(N123), .B(n77), .Z(n3) );
  CAOR2X2 U5110 ( .A(N5141), .B(n82), .C(N5237), .D(n83), .Z(N4527) );
  CAOR2X2 U5111 ( .A(N5149), .B(n82), .C(N5245), .D(n83), .Z(N3959) );
  CAOR2X2 U5112 ( .A(N5145), .B(n82), .C(N5241), .D(n83), .Z(N4243) );
  CAOR2X2 U5113 ( .A(N5138), .B(n82), .C(N5234), .D(n83), .Z(N4740) );
  CAOR2X2 U5114 ( .A(N5153), .B(n82), .C(N5249), .D(n83), .Z(N3675) );
  CAOR2X2 U5115 ( .A(N5140), .B(n82), .C(N5236), .D(n83), .Z(N4598) );
  CAOR2X2 U5116 ( .A(N5139), .B(n82), .C(N5235), .D(n83), .Z(N4669) );
  CAOR2X2 U5117 ( .A(N5143), .B(n82), .C(N5239), .D(n83), .Z(N4385) );
  CAOR2X2 U5118 ( .A(N5142), .B(n82), .C(N5238), .D(n83), .Z(N4456) );
  CAOR2X2 U5119 ( .A(N5146), .B(n82), .C(N5242), .D(n83), .Z(N4172) );
  CAOR2X2 U5120 ( .A(N5144), .B(n82), .C(N5240), .D(n83), .Z(N4314) );
  CAOR2X2 U5121 ( .A(N5148), .B(n82), .C(N5244), .D(n83), .Z(N4030) );
  CAOR2X2 U5122 ( .A(N5147), .B(n82), .C(N5243), .D(n83), .Z(N4101) );
  CAOR2X2 U5123 ( .A(N5151), .B(n82), .C(N5247), .D(n83), .Z(N3817) );
  CAOR2X2 U5124 ( .A(N5150), .B(n82), .C(N5246), .D(n83), .Z(N3888) );
  CAOR2X2 U5125 ( .A(N5154), .B(n82), .C(N5250), .D(n83), .Z(N3604) );
  CAOR2X2 U5126 ( .A(N5152), .B(n82), .C(N5248), .D(n83), .Z(N3746) );
  CAOR2X2 U5127 ( .A(N5158), .B(n82), .C(N5254), .D(n83), .Z(N3320) );
  CAOR2X2 U5128 ( .A(N5157), .B(n82), .C(N5253), .D(n83), .Z(N3391) );
  CAOR2X2 U5129 ( .A(N5156), .B(n82), .C(N5252), .D(n83), .Z(N3462) );
  CAOR2X2 U5130 ( .A(N5155), .B(n82), .C(N5251), .D(n83), .Z(N3533) );
  CAOR2X2 U5131 ( .A(N5163), .B(n82), .C(N5259), .D(n83), .Z(N2965) );
  CAOR2X2 U5132 ( .A(N5162), .B(n82), .C(N5258), .D(n83), .Z(N3036) );
  CAOR2X2 U5133 ( .A(N5160), .B(n82), .C(N5256), .D(n83), .Z(N3178) );
  CAOR2X2 U5134 ( .A(N5159), .B(n82), .C(N5255), .D(n83), .Z(N3249) );
  CIVXL U5135 ( .A(N2681), .Z(n2600) );
  CIVX2 U5136 ( .A(n2600), .Z(n2601) );
  CIVXL U5137 ( .A(N2752), .Z(n2602) );
  CIVX2 U5138 ( .A(n2602), .Z(n2603) );
  CAOR2XL U5139 ( .A(N5167), .B(n82), .C(N5263), .D(n83), .Z(N2681) );
  CAOR2XL U5140 ( .A(N5166), .B(n82), .C(N5262), .D(n83), .Z(N2752) );
  CAOR2X2 U5141 ( .A(N5165), .B(n82), .C(N5261), .D(n83), .Z(N2823) );
  CAOR2X2 U5142 ( .A(N5164), .B(n82), .C(N5260), .D(n83), .Z(N2894) );
  CIVXL U5143 ( .A(N2610), .Z(n2604) );
  CIVX2 U5144 ( .A(n2604), .Z(n2605) );
  CIVX3 U5145 ( .A(rst), .Z(n77) );
  CAOR2XL U5146 ( .A(N5168), .B(n82), .C(N5264), .D(n83), .Z(N2610) );
  CND2IXL U5147 ( .B(counter[4]), .A(counter[5]), .Z(N5107) );
  CNR2IX2 U5148 ( .B(N114), .A(N210), .Z(n2610) );
  CIVX8 U5149 ( .A(n2610), .Z(n81) );
  CIVX4 U5150 ( .A(N210), .Z(N4961) );
  COND3XL U5151 ( .A(n84), .B(N5106), .C(n85), .D(n86), .Z(N2538) );
  CAOR2X2 U5152 ( .A(N5161), .B(n82), .C(N5257), .D(n83), .Z(N3107) );
  CEOXL U5153 ( .A(counter[5]), .B(n2939), .Z(N247) );
  CEOXL U5154 ( .A(\add_116/carry[5] ), .B(counter[5]), .Z(N235) );
  COR2XL U5155 ( .A(counter[4]), .B(counter[5]), .Z(N5113) );
  CANR2XL U5156 ( .A(counter[4]), .B(n90), .C(N246), .D(n87), .Z(n88) );
  CND2XL U5157 ( .A(N4961), .B(n81), .Z(n100) );
  CEOXL U5158 ( .A(counter[4]), .B(n2938), .Z(N246) );
  CNR2IXL U5159 ( .B(n2938), .A(counter[4]), .Z(n2939) );
  CNR2X4 U5160 ( .A(N4961), .B(rst), .Z(n82) );
  CNR2X4 U5161 ( .A(n81), .B(rst), .Z(n83) );
  CAOR2X2 U5162 ( .A(N5137), .B(n82), .C(N5233), .D(n83), .Z(N4811) );
  CMX4XL U5163 ( .A0(n2929), .A1(n2927), .A2(n2928), .A3(n2926), .S0(N42), 
        .S1(N41), .Z(N44) );
  CNR2IX4 U5164 ( .B(N2539), .A(rst), .Z(N4960) );
  COR2XL U5165 ( .A(N210), .B(N4965), .Z(N2539) );
  COAN1X2 U5166 ( .A(pushin), .B(lastin), .C(N124), .Z(N5105) );
  CIVX2 U5167 ( .A(pushin), .Z(n78) );
  CIVDXL U5168 ( .A(lastin), .Z0(n79) );
  CDLY2X2 U5169 ( .A(N40), .Z(n2612) );
  CDLY2X2 U5170 ( .A(N40), .Z(n2613) );
  CDLY2X2 U5171 ( .A(N40), .Z(n2614) );
  CDLY2X2 U5172 ( .A(N40), .Z(n2615) );
  CDLY2X2 U5173 ( .A(N40), .Z(n2616) );
  CDLY2X2 U5174 ( .A(N40), .Z(n2617) );
  CDLY2X2 U5175 ( .A(N40), .Z(n2618) );
  CDLY2X2 U5176 ( .A(N40), .Z(n2619) );
  CDLY2X2 U5177 ( .A(N40), .Z(n2620) );
  CDLY2X2 U5178 ( .A(N40), .Z(n2621) );
  CDLY2X2 U5179 ( .A(N40), .Z(n2622) );
  CDLY2X2 U5180 ( .A(N40), .Z(n2623) );
  CDLY2X2 U5181 ( .A(N39), .Z(n2624) );
  CDLY2X2 U5182 ( .A(N39), .Z(n2625) );
  CDLY2X2 U5183 ( .A(N39), .Z(n2626) );
  CDLY2X2 U5184 ( .A(N39), .Z(n2627) );
  CDLY2X2 U5185 ( .A(N39), .Z(n2628) );
  CDLY2X2 U5186 ( .A(N39), .Z(n2629) );
  CDLY2X2 U5187 ( .A(N39), .Z(n2630) );
  CDLY2X2 U5188 ( .A(N39), .Z(n2631) );
  CDLY2X2 U5189 ( .A(N39), .Z(n2632) );
  CDLY2X2 U5190 ( .A(N39), .Z(n2633) );
  CDLY2X2 U5191 ( .A(N39), .Z(n2634) );
  CDLY2X2 U5192 ( .A(N39), .Z(n2635) );
  CIVXL U5193 ( .A(n2648), .Z(n2636) );
  CIVXL U5194 ( .A(n2648), .Z(n2637) );
  CIVXL U5195 ( .A(n2648), .Z(n2638) );
  CIVXL U5196 ( .A(n2648), .Z(n2639) );
  CIVXL U5197 ( .A(n2648), .Z(n2640) );
  CIVXL U5198 ( .A(n2649), .Z(n2641) );
  CIVXL U5199 ( .A(n2649), .Z(n2642) );
  CIVXL U5200 ( .A(n2649), .Z(n2643) );
  CIVXL U5201 ( .A(n2649), .Z(n2644) );
  CIVXL U5202 ( .A(n2649), .Z(n2645) );
  CIVXL U5203 ( .A(n2649), .Z(n2646) );
  CIVXL U5204 ( .A(n2649), .Z(n2647) );
  CIVX1 U5205 ( .A(N38), .Z(n2648) );
  CIVX1 U5206 ( .A(N38), .Z(n2649) );
  CMX8X1 U5207 ( .A0(\memory[24][0] ), .A1(\memory[28][0] ), .A2(
        \memory[26][0] ), .A3(\memory[30][0] ), .A4(\memory[25][0] ), .A5(
        \memory[29][0] ), .A6(\memory[27][0] ), .A7(\memory[31][0] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2650) );
  CMX8X1 U5208 ( .A0(\memory[16][0] ), .A1(\memory[20][0] ), .A2(
        \memory[18][0] ), .A3(\memory[22][0] ), .A4(\memory[17][0] ), .A5(
        \memory[21][0] ), .A6(\memory[19][0] ), .A7(\memory[23][0] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2651) );
  CMX8X1 U5209 ( .A0(\memory[8][0] ), .A1(\memory[12][0] ), .A2(
        \memory[10][0] ), .A3(\memory[14][0] ), .A4(\memory[9][0] ), .A5(
        \memory[13][0] ), .A6(\memory[11][0] ), .A7(\memory[15][0] ), .S0(
        n2617), .S1(n2629), .S2(n2642), .Z(n2652) );
  CMX8X1 U5210 ( .A0(\memory[0][0] ), .A1(\memory[4][0] ), .A2(\memory[2][0] ), 
        .A3(\memory[6][0] ), .A4(\memory[1][0] ), .A5(\memory[5][0] ), .A6(
        \memory[3][0] ), .A7(\memory[7][0] ), .S0(n2617), .S1(n2629), .S2(
        n2642), .Z(n2653) );
  CMX4X1 U5211 ( .A0(n2653), .A1(n2651), .A2(n2652), .A3(n2650), .S0(N42), 
        .S1(N41), .Z(N113) );
  CMX8X1 U5212 ( .A0(\memory[24][1] ), .A1(\memory[28][1] ), .A2(
        \memory[26][1] ), .A3(\memory[30][1] ), .A4(\memory[25][1] ), .A5(
        \memory[29][1] ), .A6(\memory[27][1] ), .A7(\memory[31][1] ), .S0(
        n2617), .S1(n2629), .S2(n2642), .Z(n2654) );
  CMX8X1 U5213 ( .A0(\memory[16][1] ), .A1(\memory[20][1] ), .A2(
        \memory[18][1] ), .A3(\memory[22][1] ), .A4(\memory[17][1] ), .A5(
        \memory[21][1] ), .A6(\memory[19][1] ), .A7(\memory[23][1] ), .S0(
        n2617), .S1(n2629), .S2(n2642), .Z(n2655) );
  CMX8X1 U5214 ( .A0(\memory[8][1] ), .A1(\memory[12][1] ), .A2(
        \memory[10][1] ), .A3(\memory[14][1] ), .A4(\memory[9][1] ), .A5(
        \memory[13][1] ), .A6(\memory[11][1] ), .A7(\memory[15][1] ), .S0(
        n2617), .S1(n2629), .S2(n2642), .Z(n2656) );
  CMX8X1 U5215 ( .A0(\memory[0][1] ), .A1(\memory[4][1] ), .A2(\memory[2][1] ), 
        .A3(\memory[6][1] ), .A4(\memory[1][1] ), .A5(\memory[5][1] ), .A6(
        \memory[3][1] ), .A7(\memory[7][1] ), .S0(n2618), .S1(n2630), .S2(
        n2642), .Z(n2657) );
  CMX4X1 U5216 ( .A0(n2657), .A1(n2655), .A2(n2656), .A3(n2654), .S0(N42), 
        .S1(N41), .Z(N112) );
  CMX8X1 U5217 ( .A0(\memory[24][2] ), .A1(\memory[28][2] ), .A2(
        \memory[26][2] ), .A3(\memory[30][2] ), .A4(\memory[25][2] ), .A5(
        \memory[29][2] ), .A6(\memory[27][2] ), .A7(\memory[31][2] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2658) );
  CMX8X1 U5218 ( .A0(\memory[16][2] ), .A1(\memory[20][2] ), .A2(
        \memory[18][2] ), .A3(\memory[22][2] ), .A4(\memory[17][2] ), .A5(
        \memory[21][2] ), .A6(\memory[19][2] ), .A7(\memory[23][2] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2659) );
  CMX8X1 U5219 ( .A0(\memory[8][2] ), .A1(\memory[12][2] ), .A2(
        \memory[10][2] ), .A3(\memory[14][2] ), .A4(\memory[9][2] ), .A5(
        \memory[13][2] ), .A6(\memory[11][2] ), .A7(\memory[15][2] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2660) );
  CMX8X1 U5220 ( .A0(\memory[0][2] ), .A1(\memory[4][2] ), .A2(\memory[2][2] ), 
        .A3(\memory[6][2] ), .A4(\memory[1][2] ), .A5(\memory[5][2] ), .A6(
        \memory[3][2] ), .A7(\memory[7][2] ), .S0(n2618), .S1(n2630), .S2(
        n2642), .Z(n2661) );
  CMX4X1 U5221 ( .A0(n2661), .A1(n2659), .A2(n2660), .A3(n2658), .S0(N42), 
        .S1(N41), .Z(N111) );
  CMX8X1 U5222 ( .A0(\memory[24][3] ), .A1(\memory[28][3] ), .A2(
        \memory[26][3] ), .A3(\memory[30][3] ), .A4(\memory[25][3] ), .A5(
        \memory[29][3] ), .A6(\memory[27][3] ), .A7(\memory[31][3] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2662) );
  CMX8X1 U5223 ( .A0(\memory[16][3] ), .A1(\memory[20][3] ), .A2(
        \memory[18][3] ), .A3(\memory[22][3] ), .A4(\memory[17][3] ), .A5(
        \memory[21][3] ), .A6(\memory[19][3] ), .A7(\memory[23][3] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2663) );
  CMX8X1 U5224 ( .A0(\memory[8][3] ), .A1(\memory[12][3] ), .A2(
        \memory[10][3] ), .A3(\memory[14][3] ), .A4(\memory[9][3] ), .A5(
        \memory[13][3] ), .A6(\memory[11][3] ), .A7(\memory[15][3] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2664) );
  CMX8X1 U5225 ( .A0(\memory[0][3] ), .A1(\memory[4][3] ), .A2(\memory[2][3] ), 
        .A3(\memory[6][3] ), .A4(\memory[1][3] ), .A5(\memory[5][3] ), .A6(
        \memory[3][3] ), .A7(\memory[7][3] ), .S0(n2618), .S1(n2630), .S2(
        n2642), .Z(n2665) );
  CMX4X1 U5226 ( .A0(n2665), .A1(n2663), .A2(n2664), .A3(n2662), .S0(N42), 
        .S1(N41), .Z(N110) );
  CMX8X1 U5227 ( .A0(\memory[24][4] ), .A1(\memory[28][4] ), .A2(
        \memory[26][4] ), .A3(\memory[30][4] ), .A4(\memory[25][4] ), .A5(
        \memory[29][4] ), .A6(\memory[27][4] ), .A7(\memory[31][4] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2666) );
  CMX8X1 U5228 ( .A0(\memory[16][4] ), .A1(\memory[20][4] ), .A2(
        \memory[18][4] ), .A3(\memory[22][4] ), .A4(\memory[17][4] ), .A5(
        \memory[21][4] ), .A6(\memory[19][4] ), .A7(\memory[23][4] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2667) );
  CMX8X1 U5229 ( .A0(\memory[8][4] ), .A1(\memory[12][4] ), .A2(
        \memory[10][4] ), .A3(\memory[14][4] ), .A4(\memory[9][4] ), .A5(
        \memory[13][4] ), .A6(\memory[11][4] ), .A7(\memory[15][4] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2668) );
  CMX8X1 U5230 ( .A0(\memory[0][4] ), .A1(\memory[4][4] ), .A2(\memory[2][4] ), 
        .A3(\memory[6][4] ), .A4(\memory[1][4] ), .A5(\memory[5][4] ), .A6(
        \memory[3][4] ), .A7(\memory[7][4] ), .S0(n2618), .S1(n2630), .S2(
        n2642), .Z(n2669) );
  CMX4X1 U5231 ( .A0(n2669), .A1(n2667), .A2(n2668), .A3(n2666), .S0(N42), 
        .S1(N41), .Z(N109) );
  CMX8X1 U5232 ( .A0(\memory[24][5] ), .A1(\memory[28][5] ), .A2(
        \memory[26][5] ), .A3(\memory[30][5] ), .A4(\memory[25][5] ), .A5(
        \memory[29][5] ), .A6(\memory[27][5] ), .A7(\memory[31][5] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2670) );
  CMX8X1 U5233 ( .A0(\memory[16][5] ), .A1(\memory[20][5] ), .A2(
        \memory[18][5] ), .A3(\memory[22][5] ), .A4(\memory[17][5] ), .A5(
        \memory[21][5] ), .A6(\memory[19][5] ), .A7(\memory[23][5] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2671) );
  CMX8X1 U5234 ( .A0(\memory[8][5] ), .A1(\memory[12][5] ), .A2(
        \memory[10][5] ), .A3(\memory[14][5] ), .A4(\memory[9][5] ), .A5(
        \memory[13][5] ), .A6(\memory[11][5] ), .A7(\memory[15][5] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2672) );
  CMX8X1 U5235 ( .A0(\memory[0][5] ), .A1(\memory[4][5] ), .A2(\memory[2][5] ), 
        .A3(\memory[6][5] ), .A4(\memory[1][5] ), .A5(\memory[5][5] ), .A6(
        \memory[3][5] ), .A7(\memory[7][5] ), .S0(n2618), .S1(n2630), .S2(
        n2642), .Z(n2673) );
  CMX4X1 U5236 ( .A0(n2673), .A1(n2671), .A2(n2672), .A3(n2670), .S0(N42), 
        .S1(N41), .Z(N108) );
  CMX8X1 U5237 ( .A0(\memory[24][6] ), .A1(\memory[28][6] ), .A2(
        \memory[26][6] ), .A3(\memory[30][6] ), .A4(\memory[25][6] ), .A5(
        \memory[29][6] ), .A6(\memory[27][6] ), .A7(\memory[31][6] ), .S0(
        n2618), .S1(n2630), .S2(n2642), .Z(n2674) );
  CMX8X1 U5238 ( .A0(\memory[16][6] ), .A1(\memory[20][6] ), .A2(
        \memory[18][6] ), .A3(\memory[22][6] ), .A4(\memory[17][6] ), .A5(
        \memory[21][6] ), .A6(\memory[19][6] ), .A7(\memory[23][6] ), .S0(
        n2618), .S1(n2630), .S2(n2643), .Z(n2675) );
  CMX8X1 U5239 ( .A0(\memory[8][6] ), .A1(\memory[12][6] ), .A2(
        \memory[10][6] ), .A3(\memory[14][6] ), .A4(\memory[9][6] ), .A5(
        \memory[13][6] ), .A6(\memory[11][6] ), .A7(\memory[15][6] ), .S0(
        n2618), .S1(n2630), .S2(n2643), .Z(n2676) );
  CMX8X1 U5240 ( .A0(\memory[0][6] ), .A1(\memory[4][6] ), .A2(\memory[2][6] ), 
        .A3(\memory[6][6] ), .A4(\memory[1][6] ), .A5(\memory[5][6] ), .A6(
        \memory[3][6] ), .A7(\memory[7][6] ), .S0(n2618), .S1(n2630), .S2(
        n2643), .Z(n2677) );
  CMX4X1 U5241 ( .A0(n2677), .A1(n2675), .A2(n2676), .A3(n2674), .S0(N42), 
        .S1(N41), .Z(N107) );
  CMX8X1 U5242 ( .A0(\memory[24][7] ), .A1(\memory[28][7] ), .A2(
        \memory[26][7] ), .A3(\memory[30][7] ), .A4(\memory[25][7] ), .A5(
        \memory[29][7] ), .A6(\memory[27][7] ), .A7(\memory[31][7] ), .S0(
        n2618), .S1(n2630), .S2(n2643), .Z(n2678) );
  CMX8X1 U5243 ( .A0(\memory[16][7] ), .A1(\memory[20][7] ), .A2(
        \memory[18][7] ), .A3(\memory[22][7] ), .A4(\memory[17][7] ), .A5(
        \memory[21][7] ), .A6(\memory[19][7] ), .A7(\memory[23][7] ), .S0(
        n2618), .S1(n2630), .S2(n2643), .Z(n2679) );
  CMX8X1 U5244 ( .A0(\memory[8][7] ), .A1(\memory[12][7] ), .A2(
        \memory[10][7] ), .A3(\memory[14][7] ), .A4(\memory[9][7] ), .A5(
        \memory[13][7] ), .A6(\memory[11][7] ), .A7(\memory[15][7] ), .S0(
        n2618), .S1(n2630), .S2(n2643), .Z(n2680) );
  CMX8X1 U5245 ( .A0(\memory[0][7] ), .A1(\memory[4][7] ), .A2(\memory[2][7] ), 
        .A3(\memory[6][7] ), .A4(\memory[1][7] ), .A5(\memory[5][7] ), .A6(
        \memory[3][7] ), .A7(\memory[7][7] ), .S0(n2618), .S1(n2630), .S2(
        n2643), .Z(n2681) );
  CMX4X1 U5246 ( .A0(n2681), .A1(n2679), .A2(n2680), .A3(n2678), .S0(N42), 
        .S1(N41), .Z(N106) );
  CMX8X1 U5247 ( .A0(\memory[24][8] ), .A1(\memory[28][8] ), .A2(
        \memory[26][8] ), .A3(\memory[30][8] ), .A4(\memory[25][8] ), .A5(
        \memory[29][8] ), .A6(\memory[27][8] ), .A7(\memory[31][8] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2682) );
  CMX8X1 U5248 ( .A0(\memory[16][8] ), .A1(\memory[20][8] ), .A2(
        \memory[18][8] ), .A3(\memory[22][8] ), .A4(\memory[17][8] ), .A5(
        \memory[21][8] ), .A6(\memory[19][8] ), .A7(\memory[23][8] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2683) );
  CMX8X1 U5249 ( .A0(\memory[8][8] ), .A1(\memory[12][8] ), .A2(
        \memory[10][8] ), .A3(\memory[14][8] ), .A4(\memory[9][8] ), .A5(
        \memory[13][8] ), .A6(\memory[11][8] ), .A7(\memory[15][8] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2684) );
  CMX8X1 U5250 ( .A0(\memory[0][8] ), .A1(\memory[4][8] ), .A2(\memory[2][8] ), 
        .A3(\memory[6][8] ), .A4(\memory[1][8] ), .A5(\memory[5][8] ), .A6(
        \memory[3][8] ), .A7(\memory[7][8] ), .S0(n2619), .S1(n2631), .S2(
        n2643), .Z(n2685) );
  CMX4X1 U5251 ( .A0(n2685), .A1(n2683), .A2(n2684), .A3(n2682), .S0(N42), 
        .S1(N41), .Z(N105) );
  CMX8X1 U5252 ( .A0(\memory[24][9] ), .A1(\memory[28][9] ), .A2(
        \memory[26][9] ), .A3(\memory[30][9] ), .A4(\memory[25][9] ), .A5(
        \memory[29][9] ), .A6(\memory[27][9] ), .A7(\memory[31][9] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2686) );
  CMX8X1 U5253 ( .A0(\memory[16][9] ), .A1(\memory[20][9] ), .A2(
        \memory[18][9] ), .A3(\memory[22][9] ), .A4(\memory[17][9] ), .A5(
        \memory[21][9] ), .A6(\memory[19][9] ), .A7(\memory[23][9] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2687) );
  CMX8X1 U5254 ( .A0(\memory[8][9] ), .A1(\memory[12][9] ), .A2(
        \memory[10][9] ), .A3(\memory[14][9] ), .A4(\memory[9][9] ), .A5(
        \memory[13][9] ), .A6(\memory[11][9] ), .A7(\memory[15][9] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2688) );
  CMX8X1 U5255 ( .A0(\memory[0][9] ), .A1(\memory[4][9] ), .A2(\memory[2][9] ), 
        .A3(\memory[6][9] ), .A4(\memory[1][9] ), .A5(\memory[5][9] ), .A6(
        \memory[3][9] ), .A7(\memory[7][9] ), .S0(n2619), .S1(n2631), .S2(
        n2643), .Z(n2689) );
  CMX4X1 U5256 ( .A0(n2689), .A1(n2687), .A2(n2688), .A3(n2686), .S0(N42), 
        .S1(N41), .Z(N104) );
  CMX8X1 U5257 ( .A0(\memory[24][10] ), .A1(\memory[28][10] ), .A2(
        \memory[26][10] ), .A3(\memory[30][10] ), .A4(\memory[25][10] ), .A5(
        \memory[29][10] ), .A6(\memory[27][10] ), .A7(\memory[31][10] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2690) );
  CMX8X1 U5258 ( .A0(\memory[16][10] ), .A1(\memory[20][10] ), .A2(
        \memory[18][10] ), .A3(\memory[22][10] ), .A4(\memory[17][10] ), .A5(
        \memory[21][10] ), .A6(\memory[19][10] ), .A7(\memory[23][10] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2691) );
  CMX8X1 U5259 ( .A0(\memory[8][10] ), .A1(\memory[12][10] ), .A2(
        \memory[10][10] ), .A3(\memory[14][10] ), .A4(\memory[9][10] ), .A5(
        \memory[13][10] ), .A6(\memory[11][10] ), .A7(\memory[15][10] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2692) );
  CMX8X1 U5260 ( .A0(\memory[0][10] ), .A1(\memory[4][10] ), .A2(
        \memory[2][10] ), .A3(\memory[6][10] ), .A4(\memory[1][10] ), .A5(
        \memory[5][10] ), .A6(\memory[3][10] ), .A7(\memory[7][10] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2693) );
  CMX4X1 U5261 ( .A0(n2693), .A1(n2691), .A2(n2692), .A3(n2690), .S0(N42), 
        .S1(N41), .Z(N103) );
  CMX8X1 U5262 ( .A0(\memory[24][11] ), .A1(\memory[28][11] ), .A2(
        \memory[26][11] ), .A3(\memory[30][11] ), .A4(\memory[25][11] ), .A5(
        \memory[29][11] ), .A6(\memory[27][11] ), .A7(\memory[31][11] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2694) );
  CMX8X1 U5263 ( .A0(\memory[16][11] ), .A1(\memory[20][11] ), .A2(
        \memory[18][11] ), .A3(\memory[22][11] ), .A4(\memory[17][11] ), .A5(
        \memory[21][11] ), .A6(\memory[19][11] ), .A7(\memory[23][11] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2695) );
  CMX8X1 U5264 ( .A0(\memory[8][11] ), .A1(\memory[12][11] ), .A2(
        \memory[10][11] ), .A3(\memory[14][11] ), .A4(\memory[9][11] ), .A5(
        \memory[13][11] ), .A6(\memory[11][11] ), .A7(\memory[15][11] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2696) );
  CMX8X1 U5265 ( .A0(\memory[0][11] ), .A1(\memory[4][11] ), .A2(
        \memory[2][11] ), .A3(\memory[6][11] ), .A4(\memory[1][11] ), .A5(
        \memory[5][11] ), .A6(\memory[3][11] ), .A7(\memory[7][11] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2697) );
  CMX4X1 U5266 ( .A0(n2697), .A1(n2695), .A2(n2696), .A3(n2694), .S0(N42), 
        .S1(N41), .Z(N102) );
  CMX8X1 U5267 ( .A0(\memory[24][12] ), .A1(\memory[28][12] ), .A2(
        \memory[26][12] ), .A3(\memory[30][12] ), .A4(\memory[25][12] ), .A5(
        \memory[29][12] ), .A6(\memory[27][12] ), .A7(\memory[31][12] ), .S0(
        n2619), .S1(n2631), .S2(n2643), .Z(n2698) );
  CMX8X1 U5268 ( .A0(\memory[16][12] ), .A1(\memory[20][12] ), .A2(
        \memory[18][12] ), .A3(\memory[22][12] ), .A4(\memory[17][12] ), .A5(
        \memory[21][12] ), .A6(\memory[19][12] ), .A7(\memory[23][12] ), .S0(
        n2619), .S1(n2631), .S2(n2644), .Z(n2699) );
  CMX8X1 U5269 ( .A0(\memory[8][12] ), .A1(\memory[12][12] ), .A2(
        \memory[10][12] ), .A3(\memory[14][12] ), .A4(\memory[9][12] ), .A5(
        \memory[13][12] ), .A6(\memory[11][12] ), .A7(\memory[15][12] ), .S0(
        n2619), .S1(n2631), .S2(n2644), .Z(n2700) );
  CMX8X1 U5270 ( .A0(\memory[0][12] ), .A1(\memory[4][12] ), .A2(
        \memory[2][12] ), .A3(\memory[6][12] ), .A4(\memory[1][12] ), .A5(
        \memory[5][12] ), .A6(\memory[3][12] ), .A7(\memory[7][12] ), .S0(
        n2619), .S1(n2631), .S2(n2644), .Z(n2701) );
  CMX4X1 U5271 ( .A0(n2701), .A1(n2699), .A2(n2700), .A3(n2698), .S0(N42), 
        .S1(N41), .Z(N101) );
  CMX8X1 U5272 ( .A0(\memory[24][13] ), .A1(\memory[28][13] ), .A2(
        \memory[26][13] ), .A3(\memory[30][13] ), .A4(\memory[25][13] ), .A5(
        \memory[29][13] ), .A6(\memory[27][13] ), .A7(\memory[31][13] ), .S0(
        n2619), .S1(n2631), .S2(n2644), .Z(n2702) );
  CMX8X1 U5273 ( .A0(\memory[16][13] ), .A1(\memory[20][13] ), .A2(
        \memory[18][13] ), .A3(\memory[22][13] ), .A4(\memory[17][13] ), .A5(
        \memory[21][13] ), .A6(\memory[19][13] ), .A7(\memory[23][13] ), .S0(
        n2619), .S1(n2631), .S2(n2644), .Z(n2703) );
  CMX8X1 U5274 ( .A0(\memory[8][13] ), .A1(\memory[12][13] ), .A2(
        \memory[10][13] ), .A3(\memory[14][13] ), .A4(\memory[9][13] ), .A5(
        \memory[13][13] ), .A6(\memory[11][13] ), .A7(\memory[15][13] ), .S0(
        n2619), .S1(n2631), .S2(n2644), .Z(n2704) );
  CMX8X1 U5275 ( .A0(\memory[0][13] ), .A1(\memory[4][13] ), .A2(
        \memory[2][13] ), .A3(\memory[6][13] ), .A4(\memory[1][13] ), .A5(
        \memory[5][13] ), .A6(\memory[3][13] ), .A7(\memory[7][13] ), .S0(
        n2619), .S1(n2631), .S2(n2644), .Z(n2705) );
  CMX4X1 U5276 ( .A0(n2705), .A1(n2703), .A2(n2704), .A3(n2702), .S0(N42), 
        .S1(N41), .Z(N100) );
  CMX8X1 U5277 ( .A0(\memory[24][14] ), .A1(\memory[28][14] ), .A2(
        \memory[26][14] ), .A3(\memory[30][14] ), .A4(\memory[25][14] ), .A5(
        \memory[29][14] ), .A6(\memory[27][14] ), .A7(\memory[31][14] ), .S0(
        n2619), .S1(n2631), .S2(n2644), .Z(n2706) );
  CMX8X1 U5278 ( .A0(\memory[16][14] ), .A1(\memory[20][14] ), .A2(
        \memory[18][14] ), .A3(\memory[22][14] ), .A4(\memory[17][14] ), .A5(
        \memory[21][14] ), .A6(\memory[19][14] ), .A7(\memory[23][14] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2707) );
  CMX8X1 U5279 ( .A0(\memory[8][14] ), .A1(\memory[12][14] ), .A2(
        \memory[10][14] ), .A3(\memory[14][14] ), .A4(\memory[9][14] ), .A5(
        \memory[13][14] ), .A6(\memory[11][14] ), .A7(\memory[15][14] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2708) );
  CMX8X1 U5280 ( .A0(\memory[0][14] ), .A1(\memory[4][14] ), .A2(
        \memory[2][14] ), .A3(\memory[6][14] ), .A4(\memory[1][14] ), .A5(
        \memory[5][14] ), .A6(\memory[3][14] ), .A7(\memory[7][14] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2709) );
  CMX4X1 U5281 ( .A0(n2709), .A1(n2707), .A2(n2708), .A3(n2706), .S0(N42), 
        .S1(N41), .Z(N99) );
  CMX8X1 U5282 ( .A0(\memory[24][15] ), .A1(\memory[28][15] ), .A2(
        \memory[26][15] ), .A3(\memory[30][15] ), .A4(\memory[25][15] ), .A5(
        \memory[29][15] ), .A6(\memory[27][15] ), .A7(\memory[31][15] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2710) );
  CMX8X1 U5283 ( .A0(\memory[16][15] ), .A1(\memory[20][15] ), .A2(
        \memory[18][15] ), .A3(\memory[22][15] ), .A4(\memory[17][15] ), .A5(
        \memory[21][15] ), .A6(\memory[19][15] ), .A7(\memory[23][15] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2711) );
  CMX8X1 U5284 ( .A0(\memory[8][15] ), .A1(\memory[12][15] ), .A2(
        \memory[10][15] ), .A3(\memory[14][15] ), .A4(\memory[9][15] ), .A5(
        \memory[13][15] ), .A6(\memory[11][15] ), .A7(\memory[15][15] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2712) );
  CMX8X1 U5285 ( .A0(\memory[0][15] ), .A1(\memory[4][15] ), .A2(
        \memory[2][15] ), .A3(\memory[6][15] ), .A4(\memory[1][15] ), .A5(
        \memory[5][15] ), .A6(\memory[3][15] ), .A7(\memory[7][15] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2713) );
  CMX4X1 U5286 ( .A0(n2713), .A1(n2711), .A2(n2712), .A3(n2710), .S0(N42), 
        .S1(N41), .Z(N98) );
  CMX8X1 U5287 ( .A0(\memory[24][16] ), .A1(\memory[28][16] ), .A2(
        \memory[26][16] ), .A3(\memory[30][16] ), .A4(\memory[25][16] ), .A5(
        \memory[29][16] ), .A6(\memory[27][16] ), .A7(\memory[31][16] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2714) );
  CMX8X1 U5288 ( .A0(\memory[16][16] ), .A1(\memory[20][16] ), .A2(
        \memory[18][16] ), .A3(\memory[22][16] ), .A4(\memory[17][16] ), .A5(
        \memory[21][16] ), .A6(\memory[19][16] ), .A7(\memory[23][16] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2715) );
  CMX8X1 U5289 ( .A0(\memory[8][16] ), .A1(\memory[12][16] ), .A2(
        \memory[10][16] ), .A3(\memory[14][16] ), .A4(\memory[9][16] ), .A5(
        \memory[13][16] ), .A6(\memory[11][16] ), .A7(\memory[15][16] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2716) );
  CMX8X1 U5290 ( .A0(\memory[0][16] ), .A1(\memory[4][16] ), .A2(
        \memory[2][16] ), .A3(\memory[6][16] ), .A4(\memory[1][16] ), .A5(
        \memory[5][16] ), .A6(\memory[3][16] ), .A7(\memory[7][16] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2717) );
  CMX4X1 U5291 ( .A0(n2717), .A1(n2715), .A2(n2716), .A3(n2714), .S0(N42), 
        .S1(N41), .Z(N97) );
  CMX8X1 U5292 ( .A0(\memory[24][17] ), .A1(\memory[28][17] ), .A2(
        \memory[26][17] ), .A3(\memory[30][17] ), .A4(\memory[25][17] ), .A5(
        \memory[29][17] ), .A6(\memory[27][17] ), .A7(\memory[31][17] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2718) );
  CMX8X1 U5293 ( .A0(\memory[16][17] ), .A1(\memory[20][17] ), .A2(
        \memory[18][17] ), .A3(\memory[22][17] ), .A4(\memory[17][17] ), .A5(
        \memory[21][17] ), .A6(\memory[19][17] ), .A7(\memory[23][17] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2719) );
  CMX8X1 U5294 ( .A0(\memory[8][17] ), .A1(\memory[12][17] ), .A2(
        \memory[10][17] ), .A3(\memory[14][17] ), .A4(\memory[9][17] ), .A5(
        \memory[13][17] ), .A6(\memory[11][17] ), .A7(\memory[15][17] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2720) );
  CMX8X1 U5295 ( .A0(\memory[0][17] ), .A1(\memory[4][17] ), .A2(
        \memory[2][17] ), .A3(\memory[6][17] ), .A4(\memory[1][17] ), .A5(
        \memory[5][17] ), .A6(\memory[3][17] ), .A7(\memory[7][17] ), .S0(
        n2620), .S1(n2632), .S2(n2644), .Z(n2721) );
  CMX4X1 U5296 ( .A0(n2721), .A1(n2719), .A2(n2720), .A3(n2718), .S0(N42), 
        .S1(N41), .Z(N96) );
  CMX8X1 U5297 ( .A0(\memory[24][18] ), .A1(\memory[28][18] ), .A2(
        \memory[26][18] ), .A3(\memory[30][18] ), .A4(\memory[25][18] ), .A5(
        \memory[29][18] ), .A6(\memory[27][18] ), .A7(\memory[31][18] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2722) );
  CMX8X1 U5298 ( .A0(\memory[16][18] ), .A1(\memory[20][18] ), .A2(
        \memory[18][18] ), .A3(\memory[22][18] ), .A4(\memory[17][18] ), .A5(
        \memory[21][18] ), .A6(\memory[19][18] ), .A7(\memory[23][18] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2723) );
  CMX8X1 U5299 ( .A0(\memory[8][18] ), .A1(\memory[12][18] ), .A2(
        \memory[10][18] ), .A3(\memory[14][18] ), .A4(\memory[9][18] ), .A5(
        \memory[13][18] ), .A6(\memory[11][18] ), .A7(\memory[15][18] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2724) );
  CMX8X1 U5300 ( .A0(\memory[0][18] ), .A1(\memory[4][18] ), .A2(
        \memory[2][18] ), .A3(\memory[6][18] ), .A4(\memory[1][18] ), .A5(
        \memory[5][18] ), .A6(\memory[3][18] ), .A7(\memory[7][18] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2725) );
  CMX4X1 U5301 ( .A0(n2725), .A1(n2723), .A2(n2724), .A3(n2722), .S0(N42), 
        .S1(N41), .Z(N95) );
  CMX8X1 U5302 ( .A0(\memory[24][19] ), .A1(\memory[28][19] ), .A2(
        \memory[26][19] ), .A3(\memory[30][19] ), .A4(\memory[25][19] ), .A5(
        \memory[29][19] ), .A6(\memory[27][19] ), .A7(\memory[31][19] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2726) );
  CMX8X1 U5303 ( .A0(\memory[16][19] ), .A1(\memory[20][19] ), .A2(
        \memory[18][19] ), .A3(\memory[22][19] ), .A4(\memory[17][19] ), .A5(
        \memory[21][19] ), .A6(\memory[19][19] ), .A7(\memory[23][19] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2727) );
  CMX8X1 U5304 ( .A0(\memory[8][19] ), .A1(\memory[12][19] ), .A2(
        \memory[10][19] ), .A3(\memory[14][19] ), .A4(\memory[9][19] ), .A5(
        \memory[13][19] ), .A6(\memory[11][19] ), .A7(\memory[15][19] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2728) );
  CMX8X1 U5305 ( .A0(\memory[0][19] ), .A1(\memory[4][19] ), .A2(
        \memory[2][19] ), .A3(\memory[6][19] ), .A4(\memory[1][19] ), .A5(
        \memory[5][19] ), .A6(\memory[3][19] ), .A7(\memory[7][19] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2729) );
  CMX4X1 U5306 ( .A0(n2729), .A1(n2727), .A2(n2728), .A3(n2726), .S0(N42), 
        .S1(N41), .Z(N94) );
  CMX8X1 U5307 ( .A0(\memory[24][20] ), .A1(\memory[28][20] ), .A2(
        \memory[26][20] ), .A3(\memory[30][20] ), .A4(\memory[25][20] ), .A5(
        \memory[29][20] ), .A6(\memory[27][20] ), .A7(\memory[31][20] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2730) );
  CMX8X1 U5308 ( .A0(\memory[16][20] ), .A1(\memory[20][20] ), .A2(
        \memory[18][20] ), .A3(\memory[22][20] ), .A4(\memory[17][20] ), .A5(
        \memory[21][20] ), .A6(\memory[19][20] ), .A7(\memory[23][20] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2731) );
  CMX8X1 U5309 ( .A0(\memory[8][20] ), .A1(\memory[12][20] ), .A2(
        \memory[10][20] ), .A3(\memory[14][20] ), .A4(\memory[9][20] ), .A5(
        \memory[13][20] ), .A6(\memory[11][20] ), .A7(\memory[15][20] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2732) );
  CMX8X1 U5310 ( .A0(\memory[0][20] ), .A1(\memory[4][20] ), .A2(
        \memory[2][20] ), .A3(\memory[6][20] ), .A4(\memory[1][20] ), .A5(
        \memory[5][20] ), .A6(\memory[3][20] ), .A7(\memory[7][20] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2733) );
  CMX4X1 U5311 ( .A0(n2733), .A1(n2731), .A2(n2732), .A3(n2730), .S0(N42), 
        .S1(N41), .Z(N93) );
  CMX8X1 U5312 ( .A0(\memory[24][21] ), .A1(\memory[28][21] ), .A2(
        \memory[26][21] ), .A3(\memory[30][21] ), .A4(\memory[25][21] ), .A5(
        \memory[29][21] ), .A6(\memory[27][21] ), .A7(\memory[31][21] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2734) );
  CMX8X1 U5313 ( .A0(\memory[16][21] ), .A1(\memory[20][21] ), .A2(
        \memory[18][21] ), .A3(\memory[22][21] ), .A4(\memory[17][21] ), .A5(
        \memory[21][21] ), .A6(\memory[19][21] ), .A7(\memory[23][21] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2735) );
  CMX8X1 U5314 ( .A0(\memory[8][21] ), .A1(\memory[12][21] ), .A2(
        \memory[10][21] ), .A3(\memory[14][21] ), .A4(\memory[9][21] ), .A5(
        \memory[13][21] ), .A6(\memory[11][21] ), .A7(\memory[15][21] ), .S0(
        n2620), .S1(n2632), .S2(n2645), .Z(n2736) );
  CMX8X1 U5315 ( .A0(\memory[0][21] ), .A1(\memory[4][21] ), .A2(
        \memory[2][21] ), .A3(\memory[6][21] ), .A4(\memory[1][21] ), .A5(
        \memory[5][21] ), .A6(\memory[3][21] ), .A7(\memory[7][21] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2737) );
  CMX4X1 U5316 ( .A0(n2737), .A1(n2735), .A2(n2736), .A3(n2734), .S0(N42), 
        .S1(N41), .Z(N92) );
  CMX8X1 U5317 ( .A0(\memory[24][22] ), .A1(\memory[28][22] ), .A2(
        \memory[26][22] ), .A3(\memory[30][22] ), .A4(\memory[25][22] ), .A5(
        \memory[29][22] ), .A6(\memory[27][22] ), .A7(\memory[31][22] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2738) );
  CMX8X1 U5318 ( .A0(\memory[16][22] ), .A1(\memory[20][22] ), .A2(
        \memory[18][22] ), .A3(\memory[22][22] ), .A4(\memory[17][22] ), .A5(
        \memory[21][22] ), .A6(\memory[19][22] ), .A7(\memory[23][22] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2739) );
  CMX8X1 U5319 ( .A0(\memory[8][22] ), .A1(\memory[12][22] ), .A2(
        \memory[10][22] ), .A3(\memory[14][22] ), .A4(\memory[9][22] ), .A5(
        \memory[13][22] ), .A6(\memory[11][22] ), .A7(\memory[15][22] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2740) );
  CMX8X1 U5320 ( .A0(\memory[0][22] ), .A1(\memory[4][22] ), .A2(
        \memory[2][22] ), .A3(\memory[6][22] ), .A4(\memory[1][22] ), .A5(
        \memory[5][22] ), .A6(\memory[3][22] ), .A7(\memory[7][22] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2741) );
  CMX4X1 U5321 ( .A0(n2741), .A1(n2739), .A2(n2740), .A3(n2738), .S0(N42), 
        .S1(N41), .Z(N91) );
  CMX8X1 U5322 ( .A0(\memory[24][23] ), .A1(\memory[28][23] ), .A2(
        \memory[26][23] ), .A3(\memory[30][23] ), .A4(\memory[25][23] ), .A5(
        \memory[29][23] ), .A6(\memory[27][23] ), .A7(\memory[31][23] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2742) );
  CMX8X1 U5323 ( .A0(\memory[16][23] ), .A1(\memory[20][23] ), .A2(
        \memory[18][23] ), .A3(\memory[22][23] ), .A4(\memory[17][23] ), .A5(
        \memory[21][23] ), .A6(\memory[19][23] ), .A7(\memory[23][23] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2743) );
  CMX8X1 U5324 ( .A0(\memory[8][23] ), .A1(\memory[12][23] ), .A2(
        \memory[10][23] ), .A3(\memory[14][23] ), .A4(\memory[9][23] ), .A5(
        \memory[13][23] ), .A6(\memory[11][23] ), .A7(\memory[15][23] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2744) );
  CMX8X1 U5325 ( .A0(\memory[0][23] ), .A1(\memory[4][23] ), .A2(
        \memory[2][23] ), .A3(\memory[6][23] ), .A4(\memory[1][23] ), .A5(
        \memory[5][23] ), .A6(\memory[3][23] ), .A7(\memory[7][23] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2745) );
  CMX4X1 U5326 ( .A0(n2745), .A1(n2743), .A2(n2744), .A3(n2742), .S0(N42), 
        .S1(N41), .Z(N90) );
  CMX8X1 U5327 ( .A0(\memory[24][24] ), .A1(\memory[28][24] ), .A2(
        \memory[26][24] ), .A3(\memory[30][24] ), .A4(\memory[25][24] ), .A5(
        \memory[29][24] ), .A6(\memory[27][24] ), .A7(\memory[31][24] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2746) );
  CMX8X1 U5328 ( .A0(\memory[16][24] ), .A1(\memory[20][24] ), .A2(
        \memory[18][24] ), .A3(\memory[22][24] ), .A4(\memory[17][24] ), .A5(
        \memory[21][24] ), .A6(\memory[19][24] ), .A7(\memory[23][24] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2747) );
  CMX8X1 U5329 ( .A0(\memory[8][24] ), .A1(\memory[12][24] ), .A2(
        \memory[10][24] ), .A3(\memory[14][24] ), .A4(\memory[9][24] ), .A5(
        \memory[13][24] ), .A6(\memory[11][24] ), .A7(\memory[15][24] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2748) );
  CMX8X1 U5330 ( .A0(\memory[0][24] ), .A1(\memory[4][24] ), .A2(
        \memory[2][24] ), .A3(\memory[6][24] ), .A4(\memory[1][24] ), .A5(
        \memory[5][24] ), .A6(\memory[3][24] ), .A7(\memory[7][24] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2749) );
  CMX4X1 U5331 ( .A0(n2749), .A1(n2747), .A2(n2748), .A3(n2746), .S0(N42), 
        .S1(N41), .Z(N89) );
  CMX8X1 U5332 ( .A0(\memory[24][25] ), .A1(\memory[28][25] ), .A2(
        \memory[26][25] ), .A3(\memory[30][25] ), .A4(\memory[25][25] ), .A5(
        \memory[29][25] ), .A6(\memory[27][25] ), .A7(\memory[31][25] ), .S0(
        n2621), .S1(n2633), .S2(n2645), .Z(n2750) );
  CMX8X1 U5333 ( .A0(\memory[16][25] ), .A1(\memory[20][25] ), .A2(
        \memory[18][25] ), .A3(\memory[22][25] ), .A4(\memory[17][25] ), .A5(
        \memory[21][25] ), .A6(\memory[19][25] ), .A7(\memory[23][25] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2751) );
  CMX8X1 U5334 ( .A0(\memory[8][25] ), .A1(\memory[12][25] ), .A2(
        \memory[10][25] ), .A3(\memory[14][25] ), .A4(\memory[9][25] ), .A5(
        \memory[13][25] ), .A6(\memory[11][25] ), .A7(\memory[15][25] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2752) );
  CMX8X1 U5335 ( .A0(\memory[0][25] ), .A1(\memory[4][25] ), .A2(
        \memory[2][25] ), .A3(\memory[6][25] ), .A4(\memory[1][25] ), .A5(
        \memory[5][25] ), .A6(\memory[3][25] ), .A7(\memory[7][25] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2753) );
  CMX4X1 U5336 ( .A0(n2753), .A1(n2751), .A2(n2752), .A3(n2750), .S0(N42), 
        .S1(N41), .Z(N88) );
  CMX8X1 U5337 ( .A0(\memory[24][26] ), .A1(\memory[28][26] ), .A2(
        \memory[26][26] ), .A3(\memory[30][26] ), .A4(\memory[25][26] ), .A5(
        \memory[29][26] ), .A6(\memory[27][26] ), .A7(\memory[31][26] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2754) );
  CMX8X1 U5338 ( .A0(\memory[16][26] ), .A1(\memory[20][26] ), .A2(
        \memory[18][26] ), .A3(\memory[22][26] ), .A4(\memory[17][26] ), .A5(
        \memory[21][26] ), .A6(\memory[19][26] ), .A7(\memory[23][26] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2755) );
  CMX8X1 U5339 ( .A0(\memory[8][26] ), .A1(\memory[12][26] ), .A2(
        \memory[10][26] ), .A3(\memory[14][26] ), .A4(\memory[9][26] ), .A5(
        \memory[13][26] ), .A6(\memory[11][26] ), .A7(\memory[15][26] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2756) );
  CMX8X1 U5340 ( .A0(\memory[0][26] ), .A1(\memory[4][26] ), .A2(
        \memory[2][26] ), .A3(\memory[6][26] ), .A4(\memory[1][26] ), .A5(
        \memory[5][26] ), .A6(\memory[3][26] ), .A7(\memory[7][26] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2757) );
  CMX4X1 U5341 ( .A0(n2757), .A1(n2755), .A2(n2756), .A3(n2754), .S0(N42), 
        .S1(N41), .Z(N87) );
  CMX8X1 U5342 ( .A0(\memory[24][27] ), .A1(\memory[28][27] ), .A2(
        \memory[26][27] ), .A3(\memory[30][27] ), .A4(\memory[25][27] ), .A5(
        \memory[29][27] ), .A6(\memory[27][27] ), .A7(\memory[31][27] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2758) );
  CMX8X1 U5343 ( .A0(\memory[16][27] ), .A1(\memory[20][27] ), .A2(
        \memory[18][27] ), .A3(\memory[22][27] ), .A4(\memory[17][27] ), .A5(
        \memory[21][27] ), .A6(\memory[19][27] ), .A7(\memory[23][27] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2759) );
  CMX8X1 U5344 ( .A0(\memory[8][27] ), .A1(\memory[12][27] ), .A2(
        \memory[10][27] ), .A3(\memory[14][27] ), .A4(\memory[9][27] ), .A5(
        \memory[13][27] ), .A6(\memory[11][27] ), .A7(\memory[15][27] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2760) );
  CMX8X1 U5345 ( .A0(\memory[0][27] ), .A1(\memory[4][27] ), .A2(
        \memory[2][27] ), .A3(\memory[6][27] ), .A4(\memory[1][27] ), .A5(
        \memory[5][27] ), .A6(\memory[3][27] ), .A7(\memory[7][27] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2761) );
  CMX4X1 U5346 ( .A0(n2761), .A1(n2759), .A2(n2760), .A3(n2758), .S0(N42), 
        .S1(N41), .Z(N86) );
  CMX8X1 U5347 ( .A0(\memory[24][28] ), .A1(\memory[28][28] ), .A2(
        \memory[26][28] ), .A3(\memory[30][28] ), .A4(\memory[25][28] ), .A5(
        \memory[29][28] ), .A6(\memory[27][28] ), .A7(\memory[31][28] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2762) );
  CMX8X1 U5348 ( .A0(\memory[16][28] ), .A1(\memory[20][28] ), .A2(
        \memory[18][28] ), .A3(\memory[22][28] ), .A4(\memory[17][28] ), .A5(
        \memory[21][28] ), .A6(\memory[19][28] ), .A7(\memory[23][28] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2763) );
  CMX8X1 U5349 ( .A0(\memory[8][28] ), .A1(\memory[12][28] ), .A2(
        \memory[10][28] ), .A3(\memory[14][28] ), .A4(\memory[9][28] ), .A5(
        \memory[13][28] ), .A6(\memory[11][28] ), .A7(\memory[15][28] ), .S0(
        n2621), .S1(n2633), .S2(n2646), .Z(n2764) );
  CMX8X1 U5350 ( .A0(\memory[0][28] ), .A1(\memory[4][28] ), .A2(
        \memory[2][28] ), .A3(\memory[6][28] ), .A4(\memory[1][28] ), .A5(
        \memory[5][28] ), .A6(\memory[3][28] ), .A7(\memory[7][28] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2765) );
  CMX4X1 U5351 ( .A0(n2765), .A1(n2763), .A2(n2764), .A3(n2762), .S0(N42), 
        .S1(N41), .Z(N85) );
  CMX8X1 U5352 ( .A0(\memory[24][29] ), .A1(\memory[28][29] ), .A2(
        \memory[26][29] ), .A3(\memory[30][29] ), .A4(\memory[25][29] ), .A5(
        \memory[29][29] ), .A6(\memory[27][29] ), .A7(\memory[31][29] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2766) );
  CMX8X1 U5353 ( .A0(\memory[16][29] ), .A1(\memory[20][29] ), .A2(
        \memory[18][29] ), .A3(\memory[22][29] ), .A4(\memory[17][29] ), .A5(
        \memory[21][29] ), .A6(\memory[19][29] ), .A7(\memory[23][29] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2767) );
  CMX8X1 U5354 ( .A0(\memory[8][29] ), .A1(\memory[12][29] ), .A2(
        \memory[10][29] ), .A3(\memory[14][29] ), .A4(\memory[9][29] ), .A5(
        \memory[13][29] ), .A6(\memory[11][29] ), .A7(\memory[15][29] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2768) );
  CMX8X1 U5355 ( .A0(\memory[0][29] ), .A1(\memory[4][29] ), .A2(
        \memory[2][29] ), .A3(\memory[6][29] ), .A4(\memory[1][29] ), .A5(
        \memory[5][29] ), .A6(\memory[3][29] ), .A7(\memory[7][29] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2769) );
  CMX4X1 U5356 ( .A0(n2769), .A1(n2767), .A2(n2768), .A3(n2766), .S0(N42), 
        .S1(N41), .Z(N84) );
  CMX8X1 U5357 ( .A0(\memory[24][30] ), .A1(\memory[28][30] ), .A2(
        \memory[26][30] ), .A3(\memory[30][30] ), .A4(\memory[25][30] ), .A5(
        \memory[29][30] ), .A6(\memory[27][30] ), .A7(\memory[31][30] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2770) );
  CMX8X1 U5358 ( .A0(\memory[16][30] ), .A1(\memory[20][30] ), .A2(
        \memory[18][30] ), .A3(\memory[22][30] ), .A4(\memory[17][30] ), .A5(
        \memory[21][30] ), .A6(\memory[19][30] ), .A7(\memory[23][30] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2771) );
  CMX8X1 U5359 ( .A0(\memory[8][30] ), .A1(\memory[12][30] ), .A2(
        \memory[10][30] ), .A3(\memory[14][30] ), .A4(\memory[9][30] ), .A5(
        \memory[13][30] ), .A6(\memory[11][30] ), .A7(\memory[15][30] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2772) );
  CMX8X1 U5360 ( .A0(\memory[0][30] ), .A1(\memory[4][30] ), .A2(
        \memory[2][30] ), .A3(\memory[6][30] ), .A4(\memory[1][30] ), .A5(
        \memory[5][30] ), .A6(\memory[3][30] ), .A7(\memory[7][30] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2773) );
  CMX4X1 U5361 ( .A0(n2773), .A1(n2771), .A2(n2772), .A3(n2770), .S0(N42), 
        .S1(N41), .Z(N83) );
  CMX8X1 U5362 ( .A0(\memory[24][31] ), .A1(\memory[28][31] ), .A2(
        \memory[26][31] ), .A3(\memory[30][31] ), .A4(\memory[25][31] ), .A5(
        \memory[29][31] ), .A6(\memory[27][31] ), .A7(\memory[31][31] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2774) );
  CMX8X1 U5363 ( .A0(\memory[16][31] ), .A1(\memory[20][31] ), .A2(
        \memory[18][31] ), .A3(\memory[22][31] ), .A4(\memory[17][31] ), .A5(
        \memory[21][31] ), .A6(\memory[19][31] ), .A7(\memory[23][31] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2775) );
  CMX8X1 U5364 ( .A0(\memory[8][31] ), .A1(\memory[12][31] ), .A2(
        \memory[10][31] ), .A3(\memory[14][31] ), .A4(\memory[9][31] ), .A5(
        \memory[13][31] ), .A6(\memory[11][31] ), .A7(\memory[15][31] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2776) );
  CMX8X1 U5365 ( .A0(\memory[0][31] ), .A1(\memory[4][31] ), .A2(
        \memory[2][31] ), .A3(\memory[6][31] ), .A4(\memory[1][31] ), .A5(
        \memory[5][31] ), .A6(\memory[3][31] ), .A7(\memory[7][31] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2777) );
  CMX4X1 U5366 ( .A0(n2777), .A1(n2775), .A2(n2776), .A3(n2774), .S0(N42), 
        .S1(N41), .Z(N82) );
  CMX8X1 U5367 ( .A0(\memory[24][32] ), .A1(\memory[28][32] ), .A2(
        \memory[26][32] ), .A3(\memory[30][32] ), .A4(\memory[25][32] ), .A5(
        \memory[29][32] ), .A6(\memory[27][32] ), .A7(\memory[31][32] ), .S0(
        n2622), .S1(n2634), .S2(n2646), .Z(n2778) );
  CMX8X1 U5368 ( .A0(\memory[16][32] ), .A1(\memory[20][32] ), .A2(
        \memory[18][32] ), .A3(\memory[22][32] ), .A4(\memory[17][32] ), .A5(
        \memory[21][32] ), .A6(\memory[19][32] ), .A7(\memory[23][32] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2779) );
  CMX8X1 U5369 ( .A0(\memory[8][32] ), .A1(\memory[12][32] ), .A2(
        \memory[10][32] ), .A3(\memory[14][32] ), .A4(\memory[9][32] ), .A5(
        \memory[13][32] ), .A6(\memory[11][32] ), .A7(\memory[15][32] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2780) );
  CMX8X1 U5370 ( .A0(\memory[0][32] ), .A1(\memory[4][32] ), .A2(
        \memory[2][32] ), .A3(\memory[6][32] ), .A4(\memory[1][32] ), .A5(
        \memory[5][32] ), .A6(\memory[3][32] ), .A7(\memory[7][32] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2781) );
  CMX4X1 U5371 ( .A0(n2781), .A1(n2779), .A2(n2780), .A3(n2778), .S0(N42), 
        .S1(N41), .Z(N81) );
  CMX8X1 U5372 ( .A0(\memory[24][33] ), .A1(\memory[28][33] ), .A2(
        \memory[26][33] ), .A3(\memory[30][33] ), .A4(\memory[25][33] ), .A5(
        \memory[29][33] ), .A6(\memory[27][33] ), .A7(\memory[31][33] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2782) );
  CMX8X1 U5373 ( .A0(\memory[16][33] ), .A1(\memory[20][33] ), .A2(
        \memory[18][33] ), .A3(\memory[22][33] ), .A4(\memory[17][33] ), .A5(
        \memory[21][33] ), .A6(\memory[19][33] ), .A7(\memory[23][33] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2783) );
  CMX8X1 U5374 ( .A0(\memory[8][33] ), .A1(\memory[12][33] ), .A2(
        \memory[10][33] ), .A3(\memory[14][33] ), .A4(\memory[9][33] ), .A5(
        \memory[13][33] ), .A6(\memory[11][33] ), .A7(\memory[15][33] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2784) );
  CMX8X1 U5375 ( .A0(\memory[0][33] ), .A1(\memory[4][33] ), .A2(
        \memory[2][33] ), .A3(\memory[6][33] ), .A4(\memory[1][33] ), .A5(
        \memory[5][33] ), .A6(\memory[3][33] ), .A7(\memory[7][33] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2785) );
  CMX4X1 U5376 ( .A0(n2785), .A1(n2783), .A2(n2784), .A3(n2782), .S0(N42), 
        .S1(N41), .Z(N80) );
  CMX8X1 U5377 ( .A0(\memory[24][34] ), .A1(\memory[28][34] ), .A2(
        \memory[26][34] ), .A3(\memory[30][34] ), .A4(\memory[25][34] ), .A5(
        \memory[29][34] ), .A6(\memory[27][34] ), .A7(\memory[31][34] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2786) );
  CMX8X1 U5378 ( .A0(\memory[16][34] ), .A1(\memory[20][34] ), .A2(
        \memory[18][34] ), .A3(\memory[22][34] ), .A4(\memory[17][34] ), .A5(
        \memory[21][34] ), .A6(\memory[19][34] ), .A7(\memory[23][34] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2787) );
  CMX8X1 U5379 ( .A0(\memory[8][34] ), .A1(\memory[12][34] ), .A2(
        \memory[10][34] ), .A3(\memory[14][34] ), .A4(\memory[9][34] ), .A5(
        \memory[13][34] ), .A6(\memory[11][34] ), .A7(\memory[15][34] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2788) );
  CMX8X1 U5380 ( .A0(\memory[0][34] ), .A1(\memory[4][34] ), .A2(
        \memory[2][34] ), .A3(\memory[6][34] ), .A4(\memory[1][34] ), .A5(
        \memory[5][34] ), .A6(\memory[3][34] ), .A7(\memory[7][34] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2789) );
  CMX4X1 U5381 ( .A0(n2789), .A1(n2787), .A2(n2788), .A3(n2786), .S0(N42), 
        .S1(N41), .Z(N79) );
  CMX8X1 U5382 ( .A0(\memory[24][35] ), .A1(\memory[28][35] ), .A2(
        \memory[26][35] ), .A3(\memory[30][35] ), .A4(\memory[25][35] ), .A5(
        \memory[29][35] ), .A6(\memory[27][35] ), .A7(\memory[31][35] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2790) );
  CMX8X1 U5383 ( .A0(\memory[16][35] ), .A1(\memory[20][35] ), .A2(
        \memory[18][35] ), .A3(\memory[22][35] ), .A4(\memory[17][35] ), .A5(
        \memory[21][35] ), .A6(\memory[19][35] ), .A7(\memory[23][35] ), .S0(
        n2623), .S1(n2635), .S2(n2647), .Z(n2791) );
  CMX8X1 U5384 ( .A0(\memory[8][35] ), .A1(\memory[12][35] ), .A2(
        \memory[10][35] ), .A3(\memory[14][35] ), .A4(\memory[9][35] ), .A5(
        \memory[13][35] ), .A6(\memory[11][35] ), .A7(\memory[15][35] ), .S0(
        n2622), .S1(n2634), .S2(n2647), .Z(n2792) );
  CMX8X1 U5385 ( .A0(\memory[0][35] ), .A1(\memory[4][35] ), .A2(
        \memory[2][35] ), .A3(\memory[6][35] ), .A4(\memory[1][35] ), .A5(
        \memory[5][35] ), .A6(\memory[3][35] ), .A7(\memory[7][35] ), .S0(
        n2614), .S1(n2626), .S2(n2639), .Z(n2793) );
  CMX4X1 U5386 ( .A0(n2793), .A1(n2791), .A2(n2792), .A3(n2790), .S0(N42), 
        .S1(N41), .Z(N78) );
  CMX8X1 U5387 ( .A0(\memory[24][36] ), .A1(\memory[28][36] ), .A2(
        \memory[26][36] ), .A3(\memory[30][36] ), .A4(\memory[25][36] ), .A5(
        \memory[29][36] ), .A6(\memory[27][36] ), .A7(\memory[31][36] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2794) );
  CMX8X1 U5388 ( .A0(\memory[16][36] ), .A1(\memory[20][36] ), .A2(
        \memory[18][36] ), .A3(\memory[22][36] ), .A4(\memory[17][36] ), .A5(
        \memory[21][36] ), .A6(\memory[19][36] ), .A7(\memory[23][36] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2795) );
  CMX8X1 U5389 ( .A0(\memory[8][36] ), .A1(\memory[12][36] ), .A2(
        \memory[10][36] ), .A3(\memory[14][36] ), .A4(\memory[9][36] ), .A5(
        \memory[13][36] ), .A6(\memory[11][36] ), .A7(\memory[15][36] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2796) );
  CMX8X1 U5390 ( .A0(\memory[0][36] ), .A1(\memory[4][36] ), .A2(
        \memory[2][36] ), .A3(\memory[6][36] ), .A4(\memory[1][36] ), .A5(
        \memory[5][36] ), .A6(\memory[3][36] ), .A7(\memory[7][36] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2797) );
  CMX4X1 U5391 ( .A0(n2797), .A1(n2795), .A2(n2796), .A3(n2794), .S0(N42), 
        .S1(N41), .Z(N77) );
  CMX8X1 U5392 ( .A0(\memory[24][37] ), .A1(\memory[28][37] ), .A2(
        \memory[26][37] ), .A3(\memory[30][37] ), .A4(\memory[25][37] ), .A5(
        \memory[29][37] ), .A6(\memory[27][37] ), .A7(\memory[31][37] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2798) );
  CMX8X1 U5393 ( .A0(\memory[16][37] ), .A1(\memory[20][37] ), .A2(
        \memory[18][37] ), .A3(\memory[22][37] ), .A4(\memory[17][37] ), .A5(
        \memory[21][37] ), .A6(\memory[19][37] ), .A7(\memory[23][37] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2799) );
  CMX8X1 U5394 ( .A0(\memory[8][37] ), .A1(\memory[12][37] ), .A2(
        \memory[10][37] ), .A3(\memory[14][37] ), .A4(\memory[9][37] ), .A5(
        \memory[13][37] ), .A6(\memory[11][37] ), .A7(\memory[15][37] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2800) );
  CMX8X1 U5395 ( .A0(\memory[0][37] ), .A1(\memory[4][37] ), .A2(
        \memory[2][37] ), .A3(\memory[6][37] ), .A4(\memory[1][37] ), .A5(
        \memory[5][37] ), .A6(\memory[3][37] ), .A7(\memory[7][37] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2801) );
  CMX4X1 U5396 ( .A0(n2801), .A1(n2799), .A2(n2800), .A3(n2798), .S0(N42), 
        .S1(N41), .Z(N76) );
  CMX8X1 U5397 ( .A0(\memory[24][38] ), .A1(\memory[28][38] ), .A2(
        \memory[26][38] ), .A3(\memory[30][38] ), .A4(\memory[25][38] ), .A5(
        \memory[29][38] ), .A6(\memory[27][38] ), .A7(\memory[31][38] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2802) );
  CMX8X1 U5398 ( .A0(\memory[16][38] ), .A1(\memory[20][38] ), .A2(
        \memory[18][38] ), .A3(\memory[22][38] ), .A4(\memory[17][38] ), .A5(
        \memory[21][38] ), .A6(\memory[19][38] ), .A7(\memory[23][38] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2803) );
  CMX8X1 U5399 ( .A0(\memory[8][38] ), .A1(\memory[12][38] ), .A2(
        \memory[10][38] ), .A3(\memory[14][38] ), .A4(\memory[9][38] ), .A5(
        \memory[13][38] ), .A6(\memory[11][38] ), .A7(\memory[15][38] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2804) );
  CMX8X1 U5400 ( .A0(\memory[0][38] ), .A1(\memory[4][38] ), .A2(
        \memory[2][38] ), .A3(\memory[6][38] ), .A4(\memory[1][38] ), .A5(
        \memory[5][38] ), .A6(\memory[3][38] ), .A7(\memory[7][38] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2805) );
  CMX4X1 U5401 ( .A0(n2805), .A1(n2803), .A2(n2804), .A3(n2802), .S0(N42), 
        .S1(N41), .Z(N75) );
  CMX8X1 U5402 ( .A0(\memory[24][39] ), .A1(\memory[28][39] ), .A2(
        \memory[26][39] ), .A3(\memory[30][39] ), .A4(\memory[25][39] ), .A5(
        \memory[29][39] ), .A6(\memory[27][39] ), .A7(\memory[31][39] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2806) );
  CMX8X1 U5403 ( .A0(\memory[16][39] ), .A1(\memory[20][39] ), .A2(
        \memory[18][39] ), .A3(\memory[22][39] ), .A4(\memory[17][39] ), .A5(
        \memory[21][39] ), .A6(\memory[19][39] ), .A7(\memory[23][39] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2807) );
  CMX8X1 U5404 ( .A0(\memory[8][39] ), .A1(\memory[12][39] ), .A2(
        \memory[10][39] ), .A3(\memory[14][39] ), .A4(\memory[9][39] ), .A5(
        \memory[13][39] ), .A6(\memory[11][39] ), .A7(\memory[15][39] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2808) );
  CMX8X1 U5405 ( .A0(\memory[0][39] ), .A1(\memory[4][39] ), .A2(
        \memory[2][39] ), .A3(\memory[6][39] ), .A4(\memory[1][39] ), .A5(
        \memory[5][39] ), .A6(\memory[3][39] ), .A7(\memory[7][39] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2809) );
  CMX4X1 U5406 ( .A0(n2809), .A1(n2807), .A2(n2808), .A3(n2806), .S0(N42), 
        .S1(N41), .Z(N74) );
  CMX8X1 U5407 ( .A0(\memory[24][40] ), .A1(\memory[28][40] ), .A2(
        \memory[26][40] ), .A3(\memory[30][40] ), .A4(\memory[25][40] ), .A5(
        \memory[29][40] ), .A6(\memory[27][40] ), .A7(\memory[31][40] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2810) );
  CMX8X1 U5408 ( .A0(\memory[16][40] ), .A1(\memory[20][40] ), .A2(
        \memory[18][40] ), .A3(\memory[22][40] ), .A4(\memory[17][40] ), .A5(
        \memory[21][40] ), .A6(\memory[19][40] ), .A7(\memory[23][40] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2811) );
  CMX8X1 U5409 ( .A0(\memory[8][40] ), .A1(\memory[12][40] ), .A2(
        \memory[10][40] ), .A3(\memory[14][40] ), .A4(\memory[9][40] ), .A5(
        \memory[13][40] ), .A6(\memory[11][40] ), .A7(\memory[15][40] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2812) );
  CMX8X1 U5410 ( .A0(\memory[0][40] ), .A1(\memory[4][40] ), .A2(
        \memory[2][40] ), .A3(\memory[6][40] ), .A4(\memory[1][40] ), .A5(
        \memory[5][40] ), .A6(\memory[3][40] ), .A7(\memory[7][40] ), .S0(
        n2612), .S1(n2624), .S2(n2636), .Z(n2813) );
  CMX4X1 U5411 ( .A0(n2813), .A1(n2811), .A2(n2812), .A3(n2810), .S0(N42), 
        .S1(N41), .Z(N73) );
  CMX8X1 U5412 ( .A0(\memory[24][41] ), .A1(\memory[28][41] ), .A2(
        \memory[26][41] ), .A3(\memory[30][41] ), .A4(\memory[25][41] ), .A5(
        \memory[29][41] ), .A6(\memory[27][41] ), .A7(\memory[31][41] ), .S0(
        n2612), .S1(n2624), .S2(n2637), .Z(n2814) );
  CMX8X1 U5413 ( .A0(\memory[16][41] ), .A1(\memory[20][41] ), .A2(
        \memory[18][41] ), .A3(\memory[22][41] ), .A4(\memory[17][41] ), .A5(
        \memory[21][41] ), .A6(\memory[19][41] ), .A7(\memory[23][41] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2815) );
  CMX8X1 U5414 ( .A0(\memory[8][41] ), .A1(\memory[12][41] ), .A2(
        \memory[10][41] ), .A3(\memory[14][41] ), .A4(\memory[9][41] ), .A5(
        \memory[13][41] ), .A6(\memory[11][41] ), .A7(\memory[15][41] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2816) );
  CMX8X1 U5415 ( .A0(\memory[0][41] ), .A1(\memory[4][41] ), .A2(
        \memory[2][41] ), .A3(\memory[6][41] ), .A4(\memory[1][41] ), .A5(
        \memory[5][41] ), .A6(\memory[3][41] ), .A7(\memory[7][41] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2817) );
  CMX4X1 U5416 ( .A0(n2817), .A1(n2815), .A2(n2816), .A3(n2814), .S0(N42), 
        .S1(N41), .Z(N72) );
  CMX8X1 U5417 ( .A0(\memory[24][42] ), .A1(\memory[28][42] ), .A2(
        \memory[26][42] ), .A3(\memory[30][42] ), .A4(\memory[25][42] ), .A5(
        \memory[29][42] ), .A6(\memory[27][42] ), .A7(\memory[31][42] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2818) );
  CMX8X1 U5418 ( .A0(\memory[16][42] ), .A1(\memory[20][42] ), .A2(
        \memory[18][42] ), .A3(\memory[22][42] ), .A4(\memory[17][42] ), .A5(
        \memory[21][42] ), .A6(\memory[19][42] ), .A7(\memory[23][42] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2819) );
  CMX8X1 U5419 ( .A0(\memory[8][42] ), .A1(\memory[12][42] ), .A2(
        \memory[10][42] ), .A3(\memory[14][42] ), .A4(\memory[9][42] ), .A5(
        \memory[13][42] ), .A6(\memory[11][42] ), .A7(\memory[15][42] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2820) );
  CMX8X1 U5420 ( .A0(\memory[0][42] ), .A1(\memory[4][42] ), .A2(
        \memory[2][42] ), .A3(\memory[6][42] ), .A4(\memory[1][42] ), .A5(
        \memory[5][42] ), .A6(\memory[3][42] ), .A7(\memory[7][42] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2821) );
  CMX4X1 U5421 ( .A0(n2821), .A1(n2819), .A2(n2820), .A3(n2818), .S0(N42), 
        .S1(N41), .Z(N71) );
  CMX8X1 U5422 ( .A0(\memory[24][43] ), .A1(\memory[28][43] ), .A2(
        \memory[26][43] ), .A3(\memory[30][43] ), .A4(\memory[25][43] ), .A5(
        \memory[29][43] ), .A6(\memory[27][43] ), .A7(\memory[31][43] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2822) );
  CMX8X1 U5423 ( .A0(\memory[16][43] ), .A1(\memory[20][43] ), .A2(
        \memory[18][43] ), .A3(\memory[22][43] ), .A4(\memory[17][43] ), .A5(
        \memory[21][43] ), .A6(\memory[19][43] ), .A7(\memory[23][43] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2823) );
  CMX8X1 U5424 ( .A0(\memory[8][43] ), .A1(\memory[12][43] ), .A2(
        \memory[10][43] ), .A3(\memory[14][43] ), .A4(\memory[9][43] ), .A5(
        \memory[13][43] ), .A6(\memory[11][43] ), .A7(\memory[15][43] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2824) );
  CMX8X1 U5425 ( .A0(\memory[0][43] ), .A1(\memory[4][43] ), .A2(
        \memory[2][43] ), .A3(\memory[6][43] ), .A4(\memory[1][43] ), .A5(
        \memory[5][43] ), .A6(\memory[3][43] ), .A7(\memory[7][43] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2825) );
  CMX4X1 U5426 ( .A0(n2825), .A1(n2823), .A2(n2824), .A3(n2822), .S0(N42), 
        .S1(N41), .Z(N70) );
  CMX8X1 U5427 ( .A0(\memory[24][44] ), .A1(\memory[28][44] ), .A2(
        \memory[26][44] ), .A3(\memory[30][44] ), .A4(\memory[25][44] ), .A5(
        \memory[29][44] ), .A6(\memory[27][44] ), .A7(\memory[31][44] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2826) );
  CMX8X1 U5428 ( .A0(\memory[16][44] ), .A1(\memory[20][44] ), .A2(
        \memory[18][44] ), .A3(\memory[22][44] ), .A4(\memory[17][44] ), .A5(
        \memory[21][44] ), .A6(\memory[19][44] ), .A7(\memory[23][44] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2827) );
  CMX8X1 U5429 ( .A0(\memory[8][44] ), .A1(\memory[12][44] ), .A2(
        \memory[10][44] ), .A3(\memory[14][44] ), .A4(\memory[9][44] ), .A5(
        \memory[13][44] ), .A6(\memory[11][44] ), .A7(\memory[15][44] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2828) );
  CMX8X1 U5430 ( .A0(\memory[0][44] ), .A1(\memory[4][44] ), .A2(
        \memory[2][44] ), .A3(\memory[6][44] ), .A4(\memory[1][44] ), .A5(
        \memory[5][44] ), .A6(\memory[3][44] ), .A7(\memory[7][44] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2829) );
  CMX4X1 U5431 ( .A0(n2829), .A1(n2827), .A2(n2828), .A3(n2826), .S0(N42), 
        .S1(N41), .Z(N69) );
  CMX8X1 U5432 ( .A0(\memory[24][45] ), .A1(\memory[28][45] ), .A2(
        \memory[26][45] ), .A3(\memory[30][45] ), .A4(\memory[25][45] ), .A5(
        \memory[29][45] ), .A6(\memory[27][45] ), .A7(\memory[31][45] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2830) );
  CMX8X1 U5433 ( .A0(\memory[16][45] ), .A1(\memory[20][45] ), .A2(
        \memory[18][45] ), .A3(\memory[22][45] ), .A4(\memory[17][45] ), .A5(
        \memory[21][45] ), .A6(\memory[19][45] ), .A7(\memory[23][45] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2831) );
  CMX8X1 U5434 ( .A0(\memory[8][45] ), .A1(\memory[12][45] ), .A2(
        \memory[10][45] ), .A3(\memory[14][45] ), .A4(\memory[9][45] ), .A5(
        \memory[13][45] ), .A6(\memory[11][45] ), .A7(\memory[15][45] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2832) );
  CMX8X1 U5435 ( .A0(\memory[0][45] ), .A1(\memory[4][45] ), .A2(
        \memory[2][45] ), .A3(\memory[6][45] ), .A4(\memory[1][45] ), .A5(
        \memory[5][45] ), .A6(\memory[3][45] ), .A7(\memory[7][45] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2833) );
  CMX4X1 U5436 ( .A0(n2833), .A1(n2831), .A2(n2832), .A3(n2830), .S0(N42), 
        .S1(N41), .Z(N68) );
  CMX8X1 U5437 ( .A0(\memory[24][46] ), .A1(\memory[28][46] ), .A2(
        \memory[26][46] ), .A3(\memory[30][46] ), .A4(\memory[25][46] ), .A5(
        \memory[29][46] ), .A6(\memory[27][46] ), .A7(\memory[31][46] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2834) );
  CMX8X1 U5438 ( .A0(\memory[16][46] ), .A1(\memory[20][46] ), .A2(
        \memory[18][46] ), .A3(\memory[22][46] ), .A4(\memory[17][46] ), .A5(
        \memory[21][46] ), .A6(\memory[19][46] ), .A7(\memory[23][46] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2835) );
  CMX8X1 U5439 ( .A0(\memory[8][46] ), .A1(\memory[12][46] ), .A2(
        \memory[10][46] ), .A3(\memory[14][46] ), .A4(\memory[9][46] ), .A5(
        \memory[13][46] ), .A6(\memory[11][46] ), .A7(\memory[15][46] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2836) );
  CMX8X1 U5440 ( .A0(\memory[0][46] ), .A1(\memory[4][46] ), .A2(
        \memory[2][46] ), .A3(\memory[6][46] ), .A4(\memory[1][46] ), .A5(
        \memory[5][46] ), .A6(\memory[3][46] ), .A7(\memory[7][46] ), .S0(
        n2613), .S1(n2625), .S2(n2637), .Z(n2837) );
  CMX4X1 U5441 ( .A0(n2837), .A1(n2835), .A2(n2836), .A3(n2834), .S0(N42), 
        .S1(N41), .Z(N67) );
  CMX8X1 U5442 ( .A0(\memory[24][47] ), .A1(\memory[28][47] ), .A2(
        \memory[26][47] ), .A3(\memory[30][47] ), .A4(\memory[25][47] ), .A5(
        \memory[29][47] ), .A6(\memory[27][47] ), .A7(\memory[31][47] ), .S0(
        n2613), .S1(n2625), .S2(n2638), .Z(n2838) );
  CMX8X1 U5443 ( .A0(\memory[16][47] ), .A1(\memory[20][47] ), .A2(
        \memory[18][47] ), .A3(\memory[22][47] ), .A4(\memory[17][47] ), .A5(
        \memory[21][47] ), .A6(\memory[19][47] ), .A7(\memory[23][47] ), .S0(
        n2613), .S1(n2625), .S2(n2638), .Z(n2839) );
  CMX8X1 U5444 ( .A0(\memory[8][47] ), .A1(\memory[12][47] ), .A2(
        \memory[10][47] ), .A3(\memory[14][47] ), .A4(\memory[9][47] ), .A5(
        \memory[13][47] ), .A6(\memory[11][47] ), .A7(\memory[15][47] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2840) );
  CMX8X1 U5445 ( .A0(\memory[0][47] ), .A1(\memory[4][47] ), .A2(
        \memory[2][47] ), .A3(\memory[6][47] ), .A4(\memory[1][47] ), .A5(
        \memory[5][47] ), .A6(\memory[3][47] ), .A7(\memory[7][47] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2841) );
  CMX4X1 U5446 ( .A0(n2841), .A1(n2839), .A2(n2840), .A3(n2838), .S0(N42), 
        .S1(N41), .Z(N66) );
  CMX8X1 U5447 ( .A0(\memory[24][48] ), .A1(\memory[28][48] ), .A2(
        \memory[26][48] ), .A3(\memory[30][48] ), .A4(\memory[25][48] ), .A5(
        \memory[29][48] ), .A6(\memory[27][48] ), .A7(\memory[31][48] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2842) );
  CMX8X1 U5448 ( .A0(\memory[16][48] ), .A1(\memory[20][48] ), .A2(
        \memory[18][48] ), .A3(\memory[22][48] ), .A4(\memory[17][48] ), .A5(
        \memory[21][48] ), .A6(\memory[19][48] ), .A7(\memory[23][48] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2843) );
  CMX8X1 U5449 ( .A0(\memory[8][48] ), .A1(\memory[12][48] ), .A2(
        \memory[10][48] ), .A3(\memory[14][48] ), .A4(\memory[9][48] ), .A5(
        \memory[13][48] ), .A6(\memory[11][48] ), .A7(\memory[15][48] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2844) );
  CMX8X1 U5450 ( .A0(\memory[0][48] ), .A1(\memory[4][48] ), .A2(
        \memory[2][48] ), .A3(\memory[6][48] ), .A4(\memory[1][48] ), .A5(
        \memory[5][48] ), .A6(\memory[3][48] ), .A7(\memory[7][48] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2845) );
  CMX4X1 U5451 ( .A0(n2845), .A1(n2843), .A2(n2844), .A3(n2842), .S0(N42), 
        .S1(N41), .Z(N65) );
  CMX8X1 U5452 ( .A0(\memory[24][49] ), .A1(\memory[28][49] ), .A2(
        \memory[26][49] ), .A3(\memory[30][49] ), .A4(\memory[25][49] ), .A5(
        \memory[29][49] ), .A6(\memory[27][49] ), .A7(\memory[31][49] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2846) );
  CMX8X1 U5453 ( .A0(\memory[16][49] ), .A1(\memory[20][49] ), .A2(
        \memory[18][49] ), .A3(\memory[22][49] ), .A4(\memory[17][49] ), .A5(
        \memory[21][49] ), .A6(\memory[19][49] ), .A7(\memory[23][49] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2847) );
  CMX8X1 U5454 ( .A0(\memory[8][49] ), .A1(\memory[12][49] ), .A2(
        \memory[10][49] ), .A3(\memory[14][49] ), .A4(\memory[9][49] ), .A5(
        \memory[13][49] ), .A6(\memory[11][49] ), .A7(\memory[15][49] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2848) );
  CMX8X1 U5455 ( .A0(\memory[0][49] ), .A1(\memory[4][49] ), .A2(
        \memory[2][49] ), .A3(\memory[6][49] ), .A4(\memory[1][49] ), .A5(
        \memory[5][49] ), .A6(\memory[3][49] ), .A7(\memory[7][49] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2849) );
  CMX4X1 U5456 ( .A0(n2849), .A1(n2847), .A2(n2848), .A3(n2846), .S0(N42), 
        .S1(N41), .Z(N64) );
  CMX8X1 U5457 ( .A0(\memory[24][50] ), .A1(\memory[28][50] ), .A2(
        \memory[26][50] ), .A3(\memory[30][50] ), .A4(\memory[25][50] ), .A5(
        \memory[29][50] ), .A6(\memory[27][50] ), .A7(\memory[31][50] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2850) );
  CMX8X1 U5458 ( .A0(\memory[16][50] ), .A1(\memory[20][50] ), .A2(
        \memory[18][50] ), .A3(\memory[22][50] ), .A4(\memory[17][50] ), .A5(
        \memory[21][50] ), .A6(\memory[19][50] ), .A7(\memory[23][50] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2851) );
  CMX8X1 U5459 ( .A0(\memory[8][50] ), .A1(\memory[12][50] ), .A2(
        \memory[10][50] ), .A3(\memory[14][50] ), .A4(\memory[9][50] ), .A5(
        \memory[13][50] ), .A6(\memory[11][50] ), .A7(\memory[15][50] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2852) );
  CMX8X1 U5460 ( .A0(\memory[0][50] ), .A1(\memory[4][50] ), .A2(
        \memory[2][50] ), .A3(\memory[6][50] ), .A4(\memory[1][50] ), .A5(
        \memory[5][50] ), .A6(\memory[3][50] ), .A7(\memory[7][50] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2853) );
  CMX4X1 U5461 ( .A0(n2853), .A1(n2851), .A2(n2852), .A3(n2850), .S0(N42), 
        .S1(N41), .Z(N63) );
  CMX8X1 U5462 ( .A0(\memory[24][51] ), .A1(\memory[28][51] ), .A2(
        \memory[26][51] ), .A3(\memory[30][51] ), .A4(\memory[25][51] ), .A5(
        \memory[29][51] ), .A6(\memory[27][51] ), .A7(\memory[31][51] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2854) );
  CMX8X1 U5463 ( .A0(\memory[16][51] ), .A1(\memory[20][51] ), .A2(
        \memory[18][51] ), .A3(\memory[22][51] ), .A4(\memory[17][51] ), .A5(
        \memory[21][51] ), .A6(\memory[19][51] ), .A7(\memory[23][51] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2855) );
  CMX8X1 U5464 ( .A0(\memory[8][51] ), .A1(\memory[12][51] ), .A2(
        \memory[10][51] ), .A3(\memory[14][51] ), .A4(\memory[9][51] ), .A5(
        \memory[13][51] ), .A6(\memory[11][51] ), .A7(\memory[15][51] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2856) );
  CMX8X1 U5465 ( .A0(\memory[0][51] ), .A1(\memory[4][51] ), .A2(
        \memory[2][51] ), .A3(\memory[6][51] ), .A4(\memory[1][51] ), .A5(
        \memory[5][51] ), .A6(\memory[3][51] ), .A7(\memory[7][51] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2857) );
  CMX4X1 U5466 ( .A0(n2857), .A1(n2855), .A2(n2856), .A3(n2854), .S0(N42), 
        .S1(N41), .Z(N62) );
  CMX8X1 U5467 ( .A0(\memory[24][52] ), .A1(\memory[28][52] ), .A2(
        \memory[26][52] ), .A3(\memory[30][52] ), .A4(\memory[25][52] ), .A5(
        \memory[29][52] ), .A6(\memory[27][52] ), .A7(\memory[31][52] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2858) );
  CMX8X1 U5468 ( .A0(\memory[16][52] ), .A1(\memory[20][52] ), .A2(
        \memory[18][52] ), .A3(\memory[22][52] ), .A4(\memory[17][52] ), .A5(
        \memory[21][52] ), .A6(\memory[19][52] ), .A7(\memory[23][52] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2859) );
  CMX8X1 U5469 ( .A0(\memory[8][52] ), .A1(\memory[12][52] ), .A2(
        \memory[10][52] ), .A3(\memory[14][52] ), .A4(\memory[9][52] ), .A5(
        \memory[13][52] ), .A6(\memory[11][52] ), .A7(\memory[15][52] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2860) );
  CMX8X1 U5470 ( .A0(\memory[0][52] ), .A1(\memory[4][52] ), .A2(
        \memory[2][52] ), .A3(\memory[6][52] ), .A4(\memory[1][52] ), .A5(
        \memory[5][52] ), .A6(\memory[3][52] ), .A7(\memory[7][52] ), .S0(
        n2614), .S1(n2626), .S2(n2638), .Z(n2861) );
  CMX4X1 U5471 ( .A0(n2861), .A1(n2859), .A2(n2860), .A3(n2858), .S0(N42), 
        .S1(N41), .Z(N61) );
  CMX8X1 U5472 ( .A0(\memory[24][53] ), .A1(\memory[28][53] ), .A2(
        \memory[26][53] ), .A3(\memory[30][53] ), .A4(\memory[25][53] ), .A5(
        \memory[29][53] ), .A6(\memory[27][53] ), .A7(\memory[31][53] ), .S0(
        n2614), .S1(n2626), .S2(n2639), .Z(n2862) );
  CMX8X1 U5473 ( .A0(\memory[16][53] ), .A1(\memory[20][53] ), .A2(
        \memory[18][53] ), .A3(\memory[22][53] ), .A4(\memory[17][53] ), .A5(
        \memory[21][53] ), .A6(\memory[19][53] ), .A7(\memory[23][53] ), .S0(
        n2614), .S1(n2626), .S2(n2639), .Z(n2863) );
  CMX8X1 U5474 ( .A0(\memory[8][53] ), .A1(\memory[12][53] ), .A2(
        \memory[10][53] ), .A3(\memory[14][53] ), .A4(\memory[9][53] ), .A5(
        \memory[13][53] ), .A6(\memory[11][53] ), .A7(\memory[15][53] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2864) );
  CMX8X1 U5475 ( .A0(\memory[0][53] ), .A1(\memory[4][53] ), .A2(
        \memory[2][53] ), .A3(\memory[6][53] ), .A4(\memory[1][53] ), .A5(
        \memory[5][53] ), .A6(\memory[3][53] ), .A7(\memory[7][53] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2865) );
  CMX4X1 U5476 ( .A0(n2865), .A1(n2863), .A2(n2864), .A3(n2862), .S0(N42), 
        .S1(N41), .Z(N60) );
  CMX8X1 U5477 ( .A0(\memory[24][54] ), .A1(\memory[28][54] ), .A2(
        \memory[26][54] ), .A3(\memory[30][54] ), .A4(\memory[25][54] ), .A5(
        \memory[29][54] ), .A6(\memory[27][54] ), .A7(\memory[31][54] ), .S0(
        n2617), .S1(n2629), .S2(n2642), .Z(n2866) );
  CMX8X1 U5478 ( .A0(\memory[16][54] ), .A1(\memory[20][54] ), .A2(
        \memory[18][54] ), .A3(\memory[22][54] ), .A4(\memory[17][54] ), .A5(
        \memory[21][54] ), .A6(\memory[19][54] ), .A7(\memory[23][54] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2867) );
  CMX8X1 U5479 ( .A0(\memory[8][54] ), .A1(\memory[12][54] ), .A2(
        \memory[10][54] ), .A3(\memory[14][54] ), .A4(\memory[9][54] ), .A5(
        \memory[13][54] ), .A6(\memory[11][54] ), .A7(\memory[15][54] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2868) );
  CMX8X1 U5480 ( .A0(\memory[0][54] ), .A1(\memory[4][54] ), .A2(
        \memory[2][54] ), .A3(\memory[6][54] ), .A4(\memory[1][54] ), .A5(
        \memory[5][54] ), .A6(\memory[3][54] ), .A7(\memory[7][54] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2869) );
  CMX4X1 U5481 ( .A0(n2869), .A1(n2867), .A2(n2868), .A3(n2866), .S0(N42), 
        .S1(N41), .Z(N59) );
  CMX8X1 U5482 ( .A0(\memory[24][55] ), .A1(\memory[28][55] ), .A2(
        \memory[26][55] ), .A3(\memory[30][55] ), .A4(\memory[25][55] ), .A5(
        \memory[29][55] ), .A6(\memory[27][55] ), .A7(\memory[31][55] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2870) );
  CMX8X1 U5483 ( .A0(\memory[16][55] ), .A1(\memory[20][55] ), .A2(
        \memory[18][55] ), .A3(\memory[22][55] ), .A4(\memory[17][55] ), .A5(
        \memory[21][55] ), .A6(\memory[19][55] ), .A7(\memory[23][55] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2871) );
  CMX8X1 U5484 ( .A0(\memory[8][55] ), .A1(\memory[12][55] ), .A2(
        \memory[10][55] ), .A3(\memory[14][55] ), .A4(\memory[9][55] ), .A5(
        \memory[13][55] ), .A6(\memory[11][55] ), .A7(\memory[15][55] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2872) );
  CMX8X1 U5485 ( .A0(\memory[0][55] ), .A1(\memory[4][55] ), .A2(
        \memory[2][55] ), .A3(\memory[6][55] ), .A4(\memory[1][55] ), .A5(
        \memory[5][55] ), .A6(\memory[3][55] ), .A7(\memory[7][55] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2873) );
  CMX4X1 U5486 ( .A0(n2873), .A1(n2871), .A2(n2872), .A3(n2870), .S0(N42), 
        .S1(N41), .Z(N58) );
  CMX8X1 U5487 ( .A0(\memory[24][56] ), .A1(\memory[28][56] ), .A2(
        \memory[26][56] ), .A3(\memory[30][56] ), .A4(\memory[25][56] ), .A5(
        \memory[29][56] ), .A6(\memory[27][56] ), .A7(\memory[31][56] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2874) );
  CMX8X1 U5488 ( .A0(\memory[16][56] ), .A1(\memory[20][56] ), .A2(
        \memory[18][56] ), .A3(\memory[22][56] ), .A4(\memory[17][56] ), .A5(
        \memory[21][56] ), .A6(\memory[19][56] ), .A7(\memory[23][56] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2875) );
  CMX8X1 U5489 ( .A0(\memory[8][56] ), .A1(\memory[12][56] ), .A2(
        \memory[10][56] ), .A3(\memory[14][56] ), .A4(\memory[9][56] ), .A5(
        \memory[13][56] ), .A6(\memory[11][56] ), .A7(\memory[15][56] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2876) );
  CMX8X1 U5490 ( .A0(\memory[0][56] ), .A1(\memory[4][56] ), .A2(
        \memory[2][56] ), .A3(\memory[6][56] ), .A4(\memory[1][56] ), .A5(
        \memory[5][56] ), .A6(\memory[3][56] ), .A7(\memory[7][56] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2877) );
  CMX4X1 U5491 ( .A0(n2877), .A1(n2875), .A2(n2876), .A3(n2874), .S0(N42), 
        .S1(N41), .Z(N57) );
  CMX8X1 U5492 ( .A0(\memory[24][57] ), .A1(\memory[28][57] ), .A2(
        \memory[26][57] ), .A3(\memory[30][57] ), .A4(\memory[25][57] ), .A5(
        \memory[29][57] ), .A6(\memory[27][57] ), .A7(\memory[31][57] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2878) );
  CMX8X1 U5493 ( .A0(\memory[16][57] ), .A1(\memory[20][57] ), .A2(
        \memory[18][57] ), .A3(\memory[22][57] ), .A4(\memory[17][57] ), .A5(
        \memory[21][57] ), .A6(\memory[19][57] ), .A7(\memory[23][57] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2879) );
  CMX8X1 U5494 ( .A0(\memory[8][57] ), .A1(\memory[12][57] ), .A2(
        \memory[10][57] ), .A3(\memory[14][57] ), .A4(\memory[9][57] ), .A5(
        \memory[13][57] ), .A6(\memory[11][57] ), .A7(\memory[15][57] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2880) );
  CMX8X1 U5495 ( .A0(\memory[0][57] ), .A1(\memory[4][57] ), .A2(
        \memory[2][57] ), .A3(\memory[6][57] ), .A4(\memory[1][57] ), .A5(
        \memory[5][57] ), .A6(\memory[3][57] ), .A7(\memory[7][57] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2881) );
  CMX4X1 U5496 ( .A0(n2881), .A1(n2879), .A2(n2880), .A3(n2878), .S0(N42), 
        .S1(N41), .Z(N56) );
  CMX8X1 U5497 ( .A0(\memory[24][58] ), .A1(\memory[28][58] ), .A2(
        \memory[26][58] ), .A3(\memory[30][58] ), .A4(\memory[25][58] ), .A5(
        \memory[29][58] ), .A6(\memory[27][58] ), .A7(\memory[31][58] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2882) );
  CMX8X1 U5498 ( .A0(\memory[16][58] ), .A1(\memory[20][58] ), .A2(
        \memory[18][58] ), .A3(\memory[22][58] ), .A4(\memory[17][58] ), .A5(
        \memory[21][58] ), .A6(\memory[19][58] ), .A7(\memory[23][58] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2883) );
  CMX8X1 U5499 ( .A0(\memory[8][58] ), .A1(\memory[12][58] ), .A2(
        \memory[10][58] ), .A3(\memory[14][58] ), .A4(\memory[9][58] ), .A5(
        \memory[13][58] ), .A6(\memory[11][58] ), .A7(\memory[15][58] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2884) );
  CMX8X1 U5500 ( .A0(\memory[0][58] ), .A1(\memory[4][58] ), .A2(
        \memory[2][58] ), .A3(\memory[6][58] ), .A4(\memory[1][58] ), .A5(
        \memory[5][58] ), .A6(\memory[3][58] ), .A7(\memory[7][58] ), .S0(
        n2615), .S1(n2627), .S2(n2639), .Z(n2885) );
  CMX4X1 U5501 ( .A0(n2885), .A1(n2883), .A2(n2884), .A3(n2882), .S0(N42), 
        .S1(N41), .Z(N55) );
  CMX8X1 U5502 ( .A0(\memory[24][59] ), .A1(\memory[28][59] ), .A2(
        \memory[26][59] ), .A3(\memory[30][59] ), .A4(\memory[25][59] ), .A5(
        \memory[29][59] ), .A6(\memory[27][59] ), .A7(\memory[31][59] ), .S0(
        n2615), .S1(n2627), .S2(n2640), .Z(n2886) );
  CMX8X1 U5503 ( .A0(\memory[16][59] ), .A1(\memory[20][59] ), .A2(
        \memory[18][59] ), .A3(\memory[22][59] ), .A4(\memory[17][59] ), .A5(
        \memory[21][59] ), .A6(\memory[19][59] ), .A7(\memory[23][59] ), .S0(
        n2615), .S1(n2627), .S2(n2640), .Z(n2887) );
  CMX8X1 U5504 ( .A0(\memory[8][59] ), .A1(\memory[12][59] ), .A2(
        \memory[10][59] ), .A3(\memory[14][59] ), .A4(\memory[9][59] ), .A5(
        \memory[13][59] ), .A6(\memory[11][59] ), .A7(\memory[15][59] ), .S0(
        n2615), .S1(n2627), .S2(n2640), .Z(n2888) );
  CMX8X1 U5505 ( .A0(\memory[0][59] ), .A1(\memory[4][59] ), .A2(
        \memory[2][59] ), .A3(\memory[6][59] ), .A4(\memory[1][59] ), .A5(
        \memory[5][59] ), .A6(\memory[3][59] ), .A7(\memory[7][59] ), .S0(
        n2615), .S1(n2627), .S2(n2640), .Z(n2889) );
  CMX4X1 U5506 ( .A0(n2889), .A1(n2887), .A2(n2888), .A3(n2886), .S0(N42), 
        .S1(N41), .Z(N54) );
  CMX8X1 U5507 ( .A0(\memory[24][60] ), .A1(\memory[28][60] ), .A2(
        \memory[26][60] ), .A3(\memory[30][60] ), .A4(\memory[25][60] ), .A5(
        \memory[29][60] ), .A6(\memory[27][60] ), .A7(\memory[31][60] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2890) );
  CMX8X1 U5508 ( .A0(\memory[16][60] ), .A1(\memory[20][60] ), .A2(
        \memory[18][60] ), .A3(\memory[22][60] ), .A4(\memory[17][60] ), .A5(
        \memory[21][60] ), .A6(\memory[19][60] ), .A7(\memory[23][60] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2891) );
  CMX8X1 U5509 ( .A0(\memory[8][60] ), .A1(\memory[12][60] ), .A2(
        \memory[10][60] ), .A3(\memory[14][60] ), .A4(\memory[9][60] ), .A5(
        \memory[13][60] ), .A6(\memory[11][60] ), .A7(\memory[15][60] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2892) );
  CMX8X1 U5510 ( .A0(\memory[0][60] ), .A1(\memory[4][60] ), .A2(
        \memory[2][60] ), .A3(\memory[6][60] ), .A4(\memory[1][60] ), .A5(
        \memory[5][60] ), .A6(\memory[3][60] ), .A7(\memory[7][60] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2893) );
  CMX4X1 U5511 ( .A0(n2893), .A1(n2891), .A2(n2892), .A3(n2890), .S0(N42), 
        .S1(N41), .Z(N53) );
  CMX8X1 U5512 ( .A0(\memory[24][61] ), .A1(\memory[28][61] ), .A2(
        \memory[26][61] ), .A3(\memory[30][61] ), .A4(\memory[25][61] ), .A5(
        \memory[29][61] ), .A6(\memory[27][61] ), .A7(\memory[31][61] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2894) );
  CMX8X1 U5513 ( .A0(\memory[16][61] ), .A1(\memory[20][61] ), .A2(
        \memory[18][61] ), .A3(\memory[22][61] ), .A4(\memory[17][61] ), .A5(
        \memory[21][61] ), .A6(\memory[19][61] ), .A7(\memory[23][61] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2895) );
  CMX8X1 U5514 ( .A0(\memory[8][61] ), .A1(\memory[12][61] ), .A2(
        \memory[10][61] ), .A3(\memory[14][61] ), .A4(\memory[9][61] ), .A5(
        \memory[13][61] ), .A6(\memory[11][61] ), .A7(\memory[15][61] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2896) );
  CMX8X1 U5515 ( .A0(\memory[0][61] ), .A1(\memory[4][61] ), .A2(
        \memory[2][61] ), .A3(\memory[6][61] ), .A4(\memory[1][61] ), .A5(
        \memory[5][61] ), .A6(\memory[3][61] ), .A7(\memory[7][61] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2897) );
  CMX4X1 U5516 ( .A0(n2897), .A1(n2895), .A2(n2896), .A3(n2894), .S0(N42), 
        .S1(N41), .Z(N52) );
  CMX8X1 U5517 ( .A0(\memory[24][62] ), .A1(\memory[28][62] ), .A2(
        \memory[26][62] ), .A3(\memory[30][62] ), .A4(\memory[25][62] ), .A5(
        \memory[29][62] ), .A6(\memory[27][62] ), .A7(\memory[31][62] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2898) );
  CMX8X1 U5518 ( .A0(\memory[16][62] ), .A1(\memory[20][62] ), .A2(
        \memory[18][62] ), .A3(\memory[22][62] ), .A4(\memory[17][62] ), .A5(
        \memory[21][62] ), .A6(\memory[19][62] ), .A7(\memory[23][62] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2899) );
  CMX8X1 U5519 ( .A0(\memory[8][62] ), .A1(\memory[12][62] ), .A2(
        \memory[10][62] ), .A3(\memory[14][62] ), .A4(\memory[9][62] ), .A5(
        \memory[13][62] ), .A6(\memory[11][62] ), .A7(\memory[15][62] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2900) );
  CMX8X1 U5520 ( .A0(\memory[0][62] ), .A1(\memory[4][62] ), .A2(
        \memory[2][62] ), .A3(\memory[6][62] ), .A4(\memory[1][62] ), .A5(
        \memory[5][62] ), .A6(\memory[3][62] ), .A7(\memory[7][62] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2901) );
  CMX4X1 U5521 ( .A0(n2901), .A1(n2899), .A2(n2900), .A3(n2898), .S0(N42), 
        .S1(N41), .Z(N51) );
  CMX8X1 U5522 ( .A0(\memory[24][63] ), .A1(\memory[28][63] ), .A2(
        \memory[26][63] ), .A3(\memory[30][63] ), .A4(\memory[25][63] ), .A5(
        \memory[29][63] ), .A6(\memory[27][63] ), .A7(\memory[31][63] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2902) );
  CMX8X1 U5523 ( .A0(\memory[16][63] ), .A1(\memory[20][63] ), .A2(
        \memory[18][63] ), .A3(\memory[22][63] ), .A4(\memory[17][63] ), .A5(
        \memory[21][63] ), .A6(\memory[19][63] ), .A7(\memory[23][63] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2903) );
  CMX8X1 U5524 ( .A0(\memory[8][63] ), .A1(\memory[12][63] ), .A2(
        \memory[10][63] ), .A3(\memory[14][63] ), .A4(\memory[9][63] ), .A5(
        \memory[13][63] ), .A6(\memory[11][63] ), .A7(\memory[15][63] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2904) );
  CMX8X1 U5525 ( .A0(\memory[0][63] ), .A1(\memory[4][63] ), .A2(
        \memory[2][63] ), .A3(\memory[6][63] ), .A4(\memory[1][63] ), .A5(
        \memory[5][63] ), .A6(\memory[3][63] ), .A7(\memory[7][63] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2905) );
  CMX4X1 U5526 ( .A0(n2905), .A1(n2903), .A2(n2904), .A3(n2902), .S0(N42), 
        .S1(N41), .Z(N50) );
  CMX8X1 U5527 ( .A0(\memory[24][64] ), .A1(\memory[28][64] ), .A2(
        \memory[26][64] ), .A3(\memory[30][64] ), .A4(\memory[25][64] ), .A5(
        \memory[29][64] ), .A6(\memory[27][64] ), .A7(\memory[31][64] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2906) );
  CMX8X1 U5528 ( .A0(\memory[16][64] ), .A1(\memory[20][64] ), .A2(
        \memory[18][64] ), .A3(\memory[22][64] ), .A4(\memory[17][64] ), .A5(
        \memory[21][64] ), .A6(\memory[19][64] ), .A7(\memory[23][64] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2907) );
  CMX8X1 U5529 ( .A0(\memory[8][64] ), .A1(\memory[12][64] ), .A2(
        \memory[10][64] ), .A3(\memory[14][64] ), .A4(\memory[9][64] ), .A5(
        \memory[13][64] ), .A6(\memory[11][64] ), .A7(\memory[15][64] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2908) );
  CMX8X1 U5530 ( .A0(\memory[0][64] ), .A1(\memory[4][64] ), .A2(
        \memory[2][64] ), .A3(\memory[6][64] ), .A4(\memory[1][64] ), .A5(
        \memory[5][64] ), .A6(\memory[3][64] ), .A7(\memory[7][64] ), .S0(
        n2616), .S1(n2628), .S2(n2640), .Z(n2909) );
  CMX4X1 U5531 ( .A0(n2909), .A1(n2907), .A2(n2908), .A3(n2906), .S0(N42), 
        .S1(N41), .Z(N49) );
  CMX8X1 U5532 ( .A0(\memory[24][65] ), .A1(\memory[28][65] ), .A2(
        \memory[26][65] ), .A3(\memory[30][65] ), .A4(\memory[25][65] ), .A5(
        \memory[29][65] ), .A6(\memory[27][65] ), .A7(\memory[31][65] ), .S0(
        n2616), .S1(n2628), .S2(n2641), .Z(n2910) );
  CMX8X1 U5533 ( .A0(\memory[16][65] ), .A1(\memory[20][65] ), .A2(
        \memory[18][65] ), .A3(\memory[22][65] ), .A4(\memory[17][65] ), .A5(
        \memory[21][65] ), .A6(\memory[19][65] ), .A7(\memory[23][65] ), .S0(
        n2616), .S1(n2628), .S2(n2641), .Z(n2911) );
  CMX8X1 U5534 ( .A0(\memory[8][65] ), .A1(\memory[12][65] ), .A2(
        \memory[10][65] ), .A3(\memory[14][65] ), .A4(\memory[9][65] ), .A5(
        \memory[13][65] ), .A6(\memory[11][65] ), .A7(\memory[15][65] ), .S0(
        n2616), .S1(n2628), .S2(n2641), .Z(n2912) );
  CMX8X1 U5535 ( .A0(\memory[0][65] ), .A1(\memory[4][65] ), .A2(
        \memory[2][65] ), .A3(\memory[6][65] ), .A4(\memory[1][65] ), .A5(
        \memory[5][65] ), .A6(\memory[3][65] ), .A7(\memory[7][65] ), .S0(
        n2616), .S1(n2628), .S2(n2641), .Z(n2913) );
  CMX4X1 U5536 ( .A0(n2913), .A1(n2911), .A2(n2912), .A3(n2910), .S0(N42), 
        .S1(N41), .Z(N48) );
  CMX8X1 U5537 ( .A0(\memory[24][66] ), .A1(\memory[28][66] ), .A2(
        \memory[26][66] ), .A3(\memory[30][66] ), .A4(\memory[25][66] ), .A5(
        \memory[29][66] ), .A6(\memory[27][66] ), .A7(\memory[31][66] ), .S0(
        n2616), .S1(n2628), .S2(n2641), .Z(n2914) );
  CMX8X1 U5538 ( .A0(\memory[16][66] ), .A1(\memory[20][66] ), .A2(
        \memory[18][66] ), .A3(\memory[22][66] ), .A4(\memory[17][66] ), .A5(
        \memory[21][66] ), .A6(\memory[19][66] ), .A7(\memory[23][66] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2915) );
  CMX8X1 U5539 ( .A0(\memory[8][66] ), .A1(\memory[12][66] ), .A2(
        \memory[10][66] ), .A3(\memory[14][66] ), .A4(\memory[9][66] ), .A5(
        \memory[13][66] ), .A6(\memory[11][66] ), .A7(\memory[15][66] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2916) );
  CMX8X1 U5540 ( .A0(\memory[0][66] ), .A1(\memory[4][66] ), .A2(
        \memory[2][66] ), .A3(\memory[6][66] ), .A4(\memory[1][66] ), .A5(
        \memory[5][66] ), .A6(\memory[3][66] ), .A7(\memory[7][66] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2917) );
  CMX4X1 U5541 ( .A0(n2917), .A1(n2915), .A2(n2916), .A3(n2914), .S0(N42), 
        .S1(N41), .Z(N47) );
  CMX8X1 U5542 ( .A0(\memory[24][67] ), .A1(\memory[28][67] ), .A2(
        \memory[26][67] ), .A3(\memory[30][67] ), .A4(\memory[25][67] ), .A5(
        \memory[29][67] ), .A6(\memory[27][67] ), .A7(\memory[31][67] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2918) );
  CMX8X1 U5543 ( .A0(\memory[16][67] ), .A1(\memory[20][67] ), .A2(
        \memory[18][67] ), .A3(\memory[22][67] ), .A4(\memory[17][67] ), .A5(
        \memory[21][67] ), .A6(\memory[19][67] ), .A7(\memory[23][67] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2919) );
  CMX8X1 U5544 ( .A0(\memory[8][67] ), .A1(\memory[12][67] ), .A2(
        \memory[10][67] ), .A3(\memory[14][67] ), .A4(\memory[9][67] ), .A5(
        \memory[13][67] ), .A6(\memory[11][67] ), .A7(\memory[15][67] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2920) );
  CMX8X1 U5545 ( .A0(\memory[0][67] ), .A1(\memory[4][67] ), .A2(
        \memory[2][67] ), .A3(\memory[6][67] ), .A4(\memory[1][67] ), .A5(
        \memory[5][67] ), .A6(\memory[3][67] ), .A7(\memory[7][67] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2921) );
  CMX4X1 U5546 ( .A0(n2921), .A1(n2919), .A2(n2920), .A3(n2918), .S0(N42), 
        .S1(N41), .Z(N46) );
  CMX8X1 U5547 ( .A0(\memory[24][68] ), .A1(\memory[28][68] ), .A2(
        \memory[26][68] ), .A3(\memory[30][68] ), .A4(\memory[25][68] ), .A5(
        \memory[29][68] ), .A6(\memory[27][68] ), .A7(\memory[31][68] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2922) );
  CMX8X1 U5548 ( .A0(\memory[16][68] ), .A1(\memory[20][68] ), .A2(
        \memory[18][68] ), .A3(\memory[22][68] ), .A4(\memory[17][68] ), .A5(
        \memory[21][68] ), .A6(\memory[19][68] ), .A7(\memory[23][68] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2923) );
  CMX8X1 U5549 ( .A0(\memory[8][68] ), .A1(\memory[12][68] ), .A2(
        \memory[10][68] ), .A3(\memory[14][68] ), .A4(\memory[9][68] ), .A5(
        \memory[13][68] ), .A6(\memory[11][68] ), .A7(\memory[15][68] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2924) );
  CMX8X1 U5550 ( .A0(\memory[0][68] ), .A1(\memory[4][68] ), .A2(
        \memory[2][68] ), .A3(\memory[6][68] ), .A4(\memory[1][68] ), .A5(
        \memory[5][68] ), .A6(\memory[3][68] ), .A7(\memory[7][68] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2925) );
  CMX4X1 U5551 ( .A0(n2925), .A1(n2923), .A2(n2924), .A3(n2922), .S0(N42), 
        .S1(N41), .Z(N45) );
  CMX8X1 U5552 ( .A0(\memory[24][69] ), .A1(\memory[28][69] ), .A2(
        \memory[26][69] ), .A3(\memory[30][69] ), .A4(\memory[25][69] ), .A5(
        \memory[29][69] ), .A6(\memory[27][69] ), .A7(\memory[31][69] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2926) );
  CMX8X1 U5553 ( .A0(\memory[16][69] ), .A1(\memory[20][69] ), .A2(
        \memory[18][69] ), .A3(\memory[22][69] ), .A4(\memory[17][69] ), .A5(
        \memory[21][69] ), .A6(\memory[19][69] ), .A7(\memory[23][69] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2927) );
  CMX8X1 U5554 ( .A0(\memory[8][69] ), .A1(\memory[12][69] ), .A2(
        \memory[10][69] ), .A3(\memory[14][69] ), .A4(\memory[9][69] ), .A5(
        \memory[13][69] ), .A6(\memory[11][69] ), .A7(\memory[15][69] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2928) );
  CMX8X1 U5555 ( .A0(\memory[0][69] ), .A1(\memory[4][69] ), .A2(
        \memory[2][69] ), .A3(\memory[6][69] ), .A4(\memory[1][69] ), .A5(
        \memory[5][69] ), .A6(\memory[3][69] ), .A7(\memory[7][69] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2929) );
  CMX8X1 U5556 ( .A0(\memory[24][70] ), .A1(\memory[28][70] ), .A2(
        \memory[26][70] ), .A3(\memory[30][70] ), .A4(\memory[25][70] ), .A5(
        \memory[29][70] ), .A6(\memory[27][70] ), .A7(\memory[31][70] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2930) );
  CMX8X1 U5557 ( .A0(\memory[16][70] ), .A1(\memory[20][70] ), .A2(
        \memory[18][70] ), .A3(\memory[22][70] ), .A4(\memory[17][70] ), .A5(
        \memory[21][70] ), .A6(\memory[19][70] ), .A7(\memory[23][70] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2931) );
  CMX8X1 U5558 ( .A0(\memory[8][70] ), .A1(\memory[12][70] ), .A2(
        \memory[10][70] ), .A3(\memory[14][70] ), .A4(\memory[9][70] ), .A5(
        \memory[13][70] ), .A6(\memory[11][70] ), .A7(\memory[15][70] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2932) );
  CMX8X1 U5559 ( .A0(\memory[0][70] ), .A1(\memory[4][70] ), .A2(
        \memory[2][70] ), .A3(\memory[6][70] ), .A4(\memory[1][70] ), .A5(
        \memory[5][70] ), .A6(\memory[3][70] ), .A7(\memory[7][70] ), .S0(
        n2617), .S1(n2629), .S2(n2641), .Z(n2933) );
  CMX4X1 U5560 ( .A0(n2933), .A1(n2931), .A2(n2932), .A3(n2930), .S0(N42), 
        .S1(N41), .Z(N43) );
  CIVX1 U5561 ( .A(write_ptr[0]), .Z(N214) );
  CEOX1 U5562 ( .A(\r183/carry[4] ), .B(write_ptr[4]), .Z(N218) );
  CEOX1 U5563 ( .A(\r184/carry[4] ), .B(N42), .Z(N223) );
  CIVX1 U5564 ( .A(counter[0]), .Z(N230) );
  CIVX1 U5565 ( .A(counter[0]), .Z(N242) );
  CNR2X1 U5566 ( .A(counter[1]), .B(counter[0]), .Z(n2934) );
  CAOR1X1 U5567 ( .A(counter[0]), .B(counter[1]), .C(n2934), .Z(N243) );
  CIVX1 U5568 ( .A(n2934), .Z(n2935) );
  CNR2X1 U5569 ( .A(n2935), .B(counter[2]), .Z(n2936) );
  CAOR1X1 U5570 ( .A(n2935), .B(counter[2]), .C(n2936), .Z(N244) );
  CIVX1 U5571 ( .A(n2936), .Z(n2937) );
  CNR2X1 U5572 ( .A(n2937), .B(counter[3]), .Z(n2938) );
  CAOR1X1 U5573 ( .A(n2937), .B(counter[3]), .C(n2938), .Z(N245) );
endmodule

